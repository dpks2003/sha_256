
//
// Verific Verilog Description of module sha_uart
//

module sha_uart (clk, rst, o_uart_tx, done);
    input clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input rst /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output o_uart_tx /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output done /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire o_uart_tx_2;
    wire n869_2;
    wire n828_2;
    wire n935_2;
    wire n940_2;
    wire n945_2;
    wire n950_2;
    wire n955_2;
    wire n868_2;
    wire n1191_2;
    
    wire \chunk_index[0] , tx_valid, \state[0] , \data_chunk[0] , n10, 
        n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, 
        n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
        n31, n32, n33, n34, n35, n36, n37, n38, n39, \useone/state[0] , 
        \useone/a[0] , \useone/b[0] , \useone/c[0] , \useone/d[0] , 
        \useone/e[0] , \useone/f[0] , \useone/g[0] , \useone/h[0] , 
        \useone/round_flag[0] , \useone/H0[0] , \useone/H1[0] , \useone/H2[0] , 
        \useone/H3[0] , \useone/H4[0] , \useone/H5[0] , \useone/H6[0] , 
        \useone/H7[0] , hashdone, \signature[0] , \useone/state[1] , 
        \useone/state[2] , \useone/a[1] , \useone/a[2] , \useone/a[3] , 
        \useone/a[4] , \useone/a[5] , \useone/a[6] , \useone/a[7] , 
        \useone/a[8] , \useone/a[9] , \useone/a[10] , \useone/a[11] , 
        \useone/a[12] , \useone/a[13] , \useone/a[14] , \useone/a[15] , 
        \useone/a[16] , \useone/a[17] , \useone/a[18] , \useone/a[19] , 
        \useone/a[20] , \useone/a[21] , \useone/a[22] , \useone/a[23] , 
        \useone/a[24] , \useone/a[25] , \useone/a[26] , \useone/a[27] , 
        \useone/a[28] , \useone/a[29] , \useone/a[30] , \useone/a[31] , 
        \useone/b[1] , \useone/b[2] , \useone/b[3] , \useone/b[4] , 
        \useone/b[5] , \useone/b[6] , \useone/b[7] , \useone/b[8] , 
        \useone/b[9] , \useone/b[10] , \useone/b[11] , \useone/b[12] , 
        \useone/b[13] , \useone/b[14] , \useone/b[15] , \useone/b[16] , 
        \useone/b[17] , \useone/b[18] , \useone/b[19] , \useone/b[20] , 
        \useone/b[21] , \useone/b[22] , \useone/b[23] , \useone/b[24] , 
        \useone/b[25] , \useone/b[26] , \useone/b[27] , \useone/b[28] , 
        \useone/b[29] , \useone/b[30] , \useone/b[31] , \useone/c[1] , 
        \useone/c[2] , \useone/c[3] , \useone/c[4] , \useone/c[5] , 
        \useone/c[6] , \useone/c[7] , \useone/c[8] , \useone/c[9] , 
        \useone/c[10] , \useone/c[11] , \useone/c[12] , \useone/c[13] , 
        \useone/c[14] , \useone/c[15] , \useone/c[16] , \useone/c[17] , 
        \useone/c[18] , \useone/c[19] , \useone/c[20] , \useone/c[21] , 
        \useone/c[22] , \useone/c[23] , \useone/c[24] , \useone/c[25] , 
        \useone/c[26] , \useone/c[27] , \useone/c[28] , \useone/c[29] , 
        \useone/c[30] , \useone/c[31] , \useone/d[1] , \useone/d[2] , 
        \useone/d[3] , \useone/d[4] , \useone/d[5] , \useone/d[6] , 
        \useone/d[7] , \useone/d[8] , \useone/d[9] , \useone/d[10] , 
        \useone/d[11] , \useone/d[12] , \useone/d[13] , \useone/d[14] , 
        \useone/d[15] , \useone/d[16] , \useone/d[17] , \useone/d[18] , 
        \useone/d[19] , \useone/d[20] , \useone/d[21] , \useone/d[22] , 
        \useone/d[23] , \useone/d[24] , \useone/d[25] , \useone/d[26] , 
        \useone/d[27] , \useone/d[28] , \useone/d[29] , \useone/d[30] , 
        \useone/d[31] , \useone/e[1] , \useone/e[2] , \useone/e[3] , 
        \useone/e[4] , \useone/e[5] , \useone/e[6] , \useone/e[7] , 
        \useone/e[8] , \useone/e[9] , \useone/e[10] , \useone/e[11] , 
        \useone/e[12] , \useone/e[13] , \useone/e[14] , \useone/e[15] , 
        \useone/e[16] , \useone/e[17] , \useone/e[18] , \useone/e[19] , 
        \useone/e[20] , \useone/e[21] , \useone/e[22] , \useone/e[23] , 
        \useone/e[24] , \useone/e[25] , \useone/e[26] , \useone/e[27] , 
        \useone/e[28] , \useone/e[29] , \useone/e[30] , \useone/e[31] , 
        \useone/f[1] , \useone/f[2] , \useone/f[3] , \useone/f[4] , 
        \useone/f[5] , \useone/f[6] , \useone/f[7] , \useone/f[8] , 
        \useone/f[9] , \useone/f[10] , \useone/f[11] , \useone/f[12] , 
        \useone/f[13] , \useone/f[14] , \useone/f[15] , \useone/f[16] , 
        \useone/f[17] , \useone/f[18] , \useone/f[19] , \useone/f[20] , 
        \useone/f[21] , \useone/f[22] , \useone/f[23] , \useone/f[24] , 
        \useone/f[25] , \useone/f[26] , \useone/f[27] , \useone/f[28] , 
        \useone/f[29] , \useone/f[30] , \useone/f[31] , \useone/g[1] , 
        \useone/g[2] , \useone/g[3] , \useone/g[4] , \useone/g[5] , 
        \useone/g[6] , \useone/g[7] , \useone/g[8] , \useone/g[9] , 
        \useone/g[10] , \useone/g[11] , \useone/g[12] , \useone/g[13] , 
        \useone/g[14] , \useone/g[15] , \useone/g[16] , \useone/g[17] , 
        \useone/g[18] , \useone/g[19] , \useone/g[20] , \useone/g[21] , 
        \useone/g[22] , \useone/g[23] , \useone/g[24] , \useone/g[25] , 
        \useone/g[26] , \useone/g[27] , \useone/g[28] , \useone/g[29] , 
        \useone/g[30] , \useone/g[31] , \useone/h[1] , \useone/h[2] , 
        \useone/h[3] , \useone/h[4] , \useone/h[5] , \useone/h[6] , 
        \useone/h[7] , \useone/h[8] , \useone/h[9] , \useone/h[10] , 
        \useone/h[11] , \useone/h[12] , \useone/h[13] , \useone/h[14] , 
        \useone/h[15] , \useone/h[16] , \useone/h[17] , \useone/h[18] , 
        \useone/h[19] , \useone/h[20] , \useone/h[21] , \useone/h[22] , 
        \useone/h[23] , \useone/h[24] , \useone/h[25] , \useone/h[26] , 
        \useone/h[27] , \useone/h[28] , \useone/h[29] , \useone/h[30] , 
        \useone/h[31] , \useone/round_flag[1] , \useone/round_flag[2] , 
        \useone/round_flag[3] , \useone/round_flag[4] , \useone/round_flag[5] , 
        \useone/round_flag[6] , \useone/H0[1] , \useone/H0[2] , \useone/H0[3] , 
        \useone/H0[4] , \useone/H0[5] , \useone/H0[6] , \useone/H0[7] , 
        \useone/H0[8] , \useone/H0[9] , \useone/H0[10] , \useone/H0[11] , 
        \useone/H0[12] , \useone/H0[13] , \useone/H0[14] , \useone/H0[15] , 
        \useone/H0[16] , \useone/H0[17] , \useone/H0[18] , \useone/H0[19] , 
        \useone/H0[20] , \useone/H0[21] , \useone/H0[22] , \useone/H0[23] , 
        \useone/H0[24] , \useone/H0[25] , \useone/H0[26] , \useone/H0[27] , 
        \useone/H0[28] , \useone/H0[29] , \useone/H0[30] , \useone/H0[31] , 
        \useone/H1[1] , \useone/H1[2] , \useone/H1[3] , \useone/H1[4] , 
        \useone/H1[5] , \useone/H1[6] , \useone/H1[7] , \useone/H1[8] , 
        \useone/H1[9] , \useone/H1[10] , \useone/H1[11] , \useone/H1[12] , 
        \useone/H1[13] , \useone/H1[14] , \useone/H1[15] , \useone/H1[16] , 
        \useone/H1[17] , \useone/H1[18] , \useone/H1[19] , \useone/H1[20] , 
        \useone/H1[21] , \useone/H1[22] , \useone/H1[23] , \useone/H1[24] , 
        \useone/H1[25] , \useone/H1[26] , \useone/H1[27] , \useone/H1[28] , 
        \useone/H1[29] , \useone/H1[30] , \useone/H1[31] , \useone/H2[1] , 
        \useone/H2[2] , \useone/H2[3] , \useone/H2[4] , \useone/H2[5] , 
        \useone/H2[6] , \useone/H2[7] , \useone/H2[8] , \useone/H2[9] , 
        \useone/H2[10] , \useone/H2[11] , \useone/H2[12] , \useone/H2[13] , 
        \useone/H2[14] , \useone/H2[15] , \useone/H2[16] , \useone/H2[17] , 
        \useone/H2[18] , \useone/H2[19] , \useone/H2[20] , \useone/H2[21] , 
        \useone/H2[22] , \useone/H2[23] , \useone/H2[24] , \useone/H2[25] , 
        \useone/H2[26] , \useone/H2[27] , \useone/H2[28] , \useone/H2[29] , 
        \useone/H2[30] , \useone/H2[31] , \useone/H3[1] , \useone/H3[2] , 
        \useone/H3[3] , \useone/H3[4] , \useone/H3[5] , \useone/H3[6] , 
        \useone/H3[7] , \useone/H3[8] , \useone/H3[9] , \useone/H3[10] , 
        \useone/H3[11] , \useone/H3[12] , \useone/H3[13] , \useone/H3[14] , 
        \useone/H3[15] , \useone/H3[16] , \useone/H3[17] , \useone/H3[18] , 
        \useone/H3[19] , \useone/H3[20] , \useone/H3[21] , \useone/H3[22] , 
        \useone/H3[23] , \useone/H3[24] , \useone/H3[25] , \useone/H3[26] , 
        \useone/H3[27] , \useone/H3[28] , \useone/H3[29] , \useone/H3[30] , 
        \useone/H3[31] , \useone/H4[1] , \useone/H4[2] , \useone/H4[3] , 
        \useone/H4[4] , \useone/H4[5] , \useone/H4[6] , \useone/H4[7] , 
        \useone/H4[8] , \useone/H4[9] , \useone/H4[10] , \useone/H4[11] , 
        \useone/H4[12] , \useone/H4[13] , \useone/H4[14] , \useone/H4[15] , 
        \useone/H4[16] , \useone/H4[17] , \useone/H4[18] , \useone/H4[19] , 
        \useone/H4[20] , \useone/H4[21] , \useone/H4[22] , \useone/H4[23] , 
        \useone/H4[24] , \useone/H4[25] , \useone/H4[26] , \useone/H4[27] , 
        \useone/H4[28] , \useone/H4[29] , \useone/H4[30] , \useone/H4[31] , 
        \useone/H5[1] , \useone/H5[2] , \useone/H5[3] , \useone/H5[4] , 
        \useone/H5[5] , \useone/H5[6] , \useone/H5[7] , \useone/H5[8] , 
        \useone/H5[9] , \useone/H5[10] , \useone/H5[11] , \useone/H5[12] , 
        \useone/H5[13] , \useone/H5[14] , \useone/H5[15] , \useone/H5[16] , 
        \useone/H5[17] , \useone/H5[18] , \useone/H5[19] , \useone/H5[20] , 
        \useone/H5[21] , \useone/H5[22] , \useone/H5[23] , \useone/H5[24] , 
        \useone/H5[25] , \useone/H5[26] , \useone/H5[27] , \useone/H5[28] , 
        \useone/H5[29] , \useone/H5[30] , \useone/H5[31] , \useone/H6[1] , 
        \useone/H6[2] , \useone/H6[3] , \useone/H6[4] , \useone/H6[5] , 
        \useone/H6[6] , \useone/H6[7] , \useone/H6[8] , \useone/H6[9] , 
        \useone/H6[10] , \useone/H6[11] , \useone/H6[12] , \useone/H6[13] , 
        \useone/H6[14] , \useone/H6[15] , \useone/H6[16] , \useone/H6[17] , 
        \useone/H6[18] , \useone/H6[19] , \useone/H6[20] , \useone/H6[21] , 
        \useone/H6[22] , \useone/H6[23] , \useone/H6[24] , \useone/H6[25] , 
        \useone/H6[26] , \useone/H6[27] , \useone/H6[28] , \useone/H6[29] , 
        \useone/H6[30] , \useone/H6[31] , \useone/H7[1] , \useone/H7[2] , 
        \useone/H7[3] , \useone/H7[4] , \useone/H7[5] , \useone/H7[6] , 
        \useone/H7[7] , \useone/H7[8] , \useone/H7[9] , \useone/H7[10] , 
        \useone/H7[11] , \useone/H7[12] , \useone/H7[13] , \useone/H7[14] , 
        \useone/H7[15] , \useone/H7[16] , \useone/H7[17] , \useone/H7[18] , 
        \useone/H7[19] , \useone/H7[20] , \useone/H7[21] , \useone/H7[22] , 
        \useone/H7[23] , \useone/H7[24] , \useone/H7[25] , \useone/H7[26] , 
        \useone/H7[27] , \useone/H7[28] , \useone/H7[29] , \useone/H7[30] , 
        \useone/H7[31] , \signature[1] , \signature[2] , \signature[3] , 
        \signature[4] , \signature[5] , \signature[6] , \signature[7] , 
        \signature[8] , \signature[9] , \signature[10] , \signature[11] , 
        \signature[12] , \signature[13] , \signature[14] , \signature[15] , 
        \signature[16] , \signature[17] , \signature[18] , \signature[19] , 
        \signature[20] , \signature[21] , \signature[22] , \signature[23] , 
        \signature[24] , \signature[25] , \signature[26] , \signature[27] , 
        \signature[28] , \signature[29] , \signature[30] , \signature[31] , 
        \signature[32] , \signature[33] , \signature[34] , \signature[35] , 
        \signature[36] , \signature[37] , \signature[38] , \signature[39] , 
        \signature[40] , \signature[41] , \signature[42] , \signature[43] , 
        \signature[44] , \signature[45] , \signature[46] , \signature[47] , 
        \signature[48] , \signature[49] , \signature[50] , \signature[51] , 
        \signature[52] , \signature[53] , \signature[54] , \signature[55] , 
        \signature[56] , \signature[57] , \signature[58] , \signature[59] , 
        \signature[60] , \signature[61] , \signature[62] , \signature[63] , 
        \signature[64] , \signature[65] , \signature[66] , \signature[67] , 
        \signature[68] , \signature[69] , \signature[70] , \signature[71] , 
        \signature[72] , \signature[73] , \signature[74] , \signature[75] , 
        \signature[76] , \signature[77] , \signature[78] , \signature[79] , 
        \signature[80] , \signature[81] , \signature[82] , \signature[83] , 
        \signature[84] , \signature[85] , \signature[86] , \signature[87] , 
        \signature[88] , \signature[89] , \signature[90] , \signature[91] , 
        \signature[92] , \signature[93] , \signature[94] , \signature[95] , 
        \signature[96] , \signature[97] , \signature[98] , \signature[99] , 
        \signature[100] , \signature[101] , \signature[102] , \signature[103] , 
        \signature[104] , \signature[105] , \signature[106] , \signature[107] , 
        \signature[108] , \signature[109] , \signature[110] , \signature[111] , 
        \signature[112] , \signature[113] , \signature[114] , \signature[115] , 
        \signature[116] , \signature[117] , \signature[118] , \signature[119] , 
        \signature[120] , \signature[121] , \signature[122] , \signature[123] , 
        \signature[124] , \signature[125] , \signature[126] , \signature[127] , 
        \signature[128] , \signature[129] , \signature[130] , \signature[131] , 
        \signature[132] , \signature[133] , \signature[134] , \signature[135] , 
        \signature[136] , \signature[137] , \signature[138] , \signature[139] , 
        \signature[140] , \signature[141] , \signature[142] , \signature[143] , 
        \signature[144] , \signature[145] , \signature[146] , \signature[147] , 
        \signature[148] , \signature[149] , \signature[150] , \signature[151] , 
        \signature[152] , \signature[153] , \signature[154] , \signature[155] , 
        \signature[156] , \signature[157] , \signature[158] , \signature[159] , 
        \signature[160] , \signature[161] , \signature[162] , \signature[163] , 
        \signature[164] , \signature[165] , \signature[166] , \signature[167] , 
        \signature[168] , \signature[169] , \signature[170] , \signature[171] , 
        \signature[172] , \signature[173] , \signature[174] , \signature[175] , 
        \signature[176] , \signature[177] , \signature[178] , \signature[179] , 
        \signature[180] , \signature[181] , \signature[182] , \signature[183] , 
        \signature[184] , \signature[185] , \signature[186] , \signature[187] , 
        \signature[188] , \signature[189] , \signature[190] , \signature[191] , 
        \signature[192] , \signature[193] , \signature[194] , \signature[195] , 
        \signature[196] , \signature[197] , \signature[198] , \signature[199] , 
        \signature[200] , \signature[201] , \signature[202] , \signature[203] , 
        \signature[204] , \signature[205] , \signature[206] , \signature[207] , 
        \signature[208] , \signature[209] , \signature[210] , \signature[211] , 
        \signature[212] , \signature[213] , \signature[214] , \signature[215] , 
        \signature[216] , \signature[217] , \signature[218] , \signature[219] , 
        \signature[220] , \signature[221] , \signature[222] , \signature[223] , 
        \signature[224] , \signature[225] , \signature[226] , \signature[227] , 
        \signature[228] , \signature[229] , \signature[230] , \signature[231] , 
        \signature[232] , \signature[233] , \signature[234] , \signature[235] , 
        \signature[236] , \signature[237] , \signature[238] , \signature[239] , 
        \signature[240] , \signature[241] , \signature[242] , \signature[243] , 
        \signature[244] , \signature[245] , \signature[246] , \signature[247] , 
        \signature[248] , \signature[249] , \signature[250] , \signature[251] , 
        \signature[252] , \signature[253] , \signature[254] , \signature[255] , 
        \useuart/r_Clock_Count[0] , \useuart/r_Bit_Index[0] , o_Tx_active, 
        \useuart/r_Tx_Data[0] , \useuart/r_SM_Main[0] , \useuart/r_Clock_Count[1] , 
        \useuart/r_Clock_Count[2] , \useuart/r_Clock_Count[3] , \useuart/r_Clock_Count[4] , 
        \useuart/r_Clock_Count[5] , \useuart/r_Clock_Count[6] , \useuart/r_Clock_Count[7] , 
        \useuart/r_Clock_Count[8] , \useuart/r_Clock_Count[9] , \useuart/r_Clock_Count[10] , 
        \useuart/r_Clock_Count[11] , \useuart/r_Clock_Count[12] , \useuart/r_Bit_Index[1] , 
        \useuart/r_Bit_Index[2] , \useuart/r_Tx_Data[1] , \useuart/r_Tx_Data[2] , 
        \useuart/r_Tx_Data[3] , \useuart/r_Tx_Data[4] , \useuart/r_Tx_Data[5] , 
        \useuart/r_Tx_Data[6] , \useuart/r_Tx_Data[7] , \chunk_index[1] , 
        \chunk_index[2] , \chunk_index[3] , \chunk_index[4] , \chunk_index[5] , 
        n861, n862, n863, n864, n865, n866, n867, n868, n869, 
        n870, n871, n872, n873, n874, n875, n876, n877, n878, 
        n879, n880, n881, n882, n883, n884, n885, n886, n887, 
        n888, n889, n890, n891, n892, n893, n894, n895, n896, 
        n897, n898, n899, n900, n901, n902, n903, n904, n905, 
        n906, n907, n908, n909, n910, n911, n912, n913, n914, 
        n915, n916, n917, n918, n919, n920, n921, n922, n923, 
        n924, n925, n926, n927, n928, n929, n930, n931, n932, 
        n933, n934, n935, n936, n937, n938, n939, n940, n941, 
        n942, n943, n944, n945, n946, n947, n948, n949, n950, 
        n951, n952, n953, n954, n955, n956, n957, n958, n959, 
        n960, n961, n962, n963, n964, n965, n966, n967, n968, 
        n969, n970, n971, n972, n973, n974, n975, n976, n977, 
        n978, n979, n980, n981, n982, n983, n984, n985, n986, 
        n987, n988, n989, n990, n991, n992, n993, n994, n995, 
        n996, n997, n998, n999, n1000, n1001, n1002, n1003, 
        n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, 
        n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
        n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
        n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
        n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
        n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, 
        n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
        n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, 
        n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, 
        n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
        n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, 
        n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
        n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
        n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, 
        n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
        n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
        n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
        n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, 
        n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, 
        n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
        n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, 
        n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
        n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, 
        n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, 
        n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
        n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, 
        n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
        n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, 
        n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, 
        n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
        n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, 
        n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
        n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, 
        n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, 
        n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
        n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, 
        n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
        n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, 
        n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, 
        n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, 
        n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, 
        n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
        n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, 
        n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
        n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, 
        n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, 
        n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
        n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, 
        n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
        n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, 
        n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, 
        n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
        n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
        n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
        n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, 
        n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, 
        n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
        n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, 
        n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
        n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, 
        n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, 
        n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
        n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, 
        n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
        n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, 
        n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, 
        n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
        n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, 
        n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
        n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, 
        n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, 
        n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
        n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, 
        n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
        n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, 
        n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, 
        n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
        n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, 
        n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
        n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, 
        n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, 
        n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
        n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, 
        n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
        n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, 
        n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, 
        n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
        n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, 
        n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
        n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
        n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, 
        n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
        n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, 
        n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, 
        n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, 
        n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, 
        n1772, n1773, n1774, n1775, \i131/useone/w[17][23] , ceg_net40, 
        ceg_net85, \state[1] , ceg_net86, ceg_net99, n1790, n1792, 
        n1794, n1796, n1797, n1798, \useone/select_1072/Select_0/n5 , 
        \useone/n144202 , \useone/select_1072/Select_2/n3 , \useone/equal_1069/n7 , 
        \useone/select_1071/Select_0/n2 , \useone/select_1072/Select_1/n8 , 
        \useone/n39302 , \useone/n46233 , \useone/n46238 , \useone/n46243 , 
        \useone/n46248 , \useone/n46253 , \useone/n46258 , \useone/select_1071/Select_1/n2 , 
        \useone/n39297 , \useone/select_1071/Select_3/n2 , \useone/select_1071/Select_4/n2 , 
        \useone/select_1071/Select_5/n2 , \useone/n39293 , \useone/select_1071/Select_7/n2 , 
        \useone/select_1071/Select_8/n2 , \useone/select_1071/Select_9/n2 , 
        \useone/select_1071/Select_10/n2 , \useone/select_1071/Select_11/n2 , 
        \useone/select_1071/Select_12/n2 , \useone/select_1071/Select_13/n2 , 
        \useone/select_1071/Select_14/n2 , \useone/n39284 , \useone/select_1071/Select_16/n2 , 
        \useone/select_1071/Select_17/n2 , \useone/select_1071/Select_18/n2 , 
        \useone/select_1071/Select_19/n2 , \useone/select_1071/Select_20/n2 , 
        \useone/select_1071/Select_21/n2 , \useone/select_1071/Select_22/n2 , 
        \useone/select_1071/Select_23/n2 , \useone/select_1071/Select_24/n2 , 
        \useone/select_1071/Select_25/n2 , \useone/select_1071/Select_26/n2 , 
        \useone/select_1071/Select_27/n2 , \useone/select_1071/Select_28/n2 , 
        \useone/select_1071/Select_29/n2 , \useone/select_1071/Select_30/n2 , 
        \useone/select_1071/Select_31/n2 , \useone/select_1071/Select_32/n2 , 
        \useone/select_1071/Select_33/n2 , \useone/select_1071/Select_34/n2 , 
        \useone/select_1071/Select_35/n2 , \useone/select_1071/Select_36/n2 , 
        \useone/select_1071/Select_37/n2 , \useone/select_1071/Select_38/n2 , 
        \useone/select_1071/Select_39/n2 , \useone/select_1071/Select_40/n2 , 
        \useone/select_1071/Select_41/n2 , \useone/select_1071/Select_42/n2 , 
        \useone/select_1071/Select_43/n2 , \useone/select_1071/Select_44/n2 , 
        \useone/select_1071/Select_45/n2 , \useone/select_1071/Select_46/n2 , 
        \useone/select_1071/Select_47/n2 , \useone/select_1071/Select_48/n2 , 
        \useone/select_1071/Select_49/n2 , \useone/select_1071/Select_50/n2 , 
        \useone/select_1071/Select_51/n2 , \useone/select_1071/Select_52/n2 , 
        \useone/select_1071/Select_53/n2 , \useone/select_1071/Select_54/n2 , 
        \useone/select_1071/Select_55/n2 , \useone/select_1071/Select_56/n2 , 
        \useone/select_1071/Select_57/n2 , \useone/select_1071/Select_58/n2 , 
        \useone/select_1071/Select_59/n2 , \useone/n39239 , \useone/select_1071/Select_61/n2 , 
        \useone/select_1071/Select_62/n2 , \useone/select_1071/Select_63/n2 , 
        \useone/select_1071/Select_64/n2 , \useone/select_1071/Select_65/n2 , 
        \useone/select_1071/Select_66/n2 , \useone/select_1071/Select_67/n2 , 
        \useone/select_1071/Select_68/n2 , \useone/select_1071/Select_69/n2 , 
        \useone/select_1071/Select_70/n2 , \useone/select_1071/Select_71/n2 , 
        \useone/select_1071/Select_72/n2 , \useone/select_1071/Select_73/n2 , 
        \useone/select_1071/Select_74/n2 , \useone/select_1071/Select_75/n2 , 
        \useone/select_1071/Select_76/n2 , \useone/select_1071/Select_77/n2 , 
        \useone/select_1071/Select_78/n2 , \useone/select_1071/Select_79/n2 , 
        \useone/select_1071/Select_80/n2 , \useone/select_1071/Select_81/n2 , 
        \useone/select_1071/Select_82/n2 , \useone/select_1071/Select_83/n2 , 
        \useone/select_1071/Select_84/n2 , \useone/select_1071/Select_85/n2 , 
        \useone/select_1071/Select_86/n2 , \useone/select_1071/Select_87/n2 , 
        \useone/select_1071/Select_88/n2 , \useone/select_1071/Select_89/n2 , 
        \useone/select_1071/Select_90/n2 , \useone/select_1071/Select_91/n2 , 
        \useone/select_1071/Select_92/n2 , \useone/select_1071/Select_93/n2 , 
        \useone/select_1071/Select_94/n2 , \useone/select_1071/Select_95/n2 , 
        \useone/select_1071/Select_96/n2 , \useone/select_1071/Select_97/n2 , 
        \useone/select_1071/Select_98/n2 , \useone/select_1071/Select_99/n2 , 
        \useone/select_1071/Select_100/n2 , \useone/select_1071/Select_101/n2 , 
        \useone/select_1071/Select_102/n2 , \useone/select_1071/Select_103/n2 , 
        \useone/select_1071/Select_104/n2 , \useone/select_1071/Select_105/n2 , 
        \useone/select_1071/Select_106/n2 , \useone/select_1071/Select_107/n2 , 
        \useone/select_1071/Select_108/n2 , \useone/select_1071/Select_109/n2 , 
        \useone/select_1071/Select_110/n2 , \useone/select_1071/Select_111/n2 , 
        \useone/select_1071/Select_112/n2 , \useone/select_1071/Select_113/n2 , 
        \useone/select_1071/Select_114/n2 , \useone/select_1071/Select_115/n2 , 
        \useone/select_1071/Select_116/n2 , \useone/select_1071/Select_117/n2 , 
        \useone/select_1071/Select_118/n2 , \useone/select_1071/Select_119/n2 , 
        \useone/select_1071/Select_120/n2 , \useone/select_1071/Select_121/n2 , 
        \useone/select_1071/Select_122/n2 , \useone/select_1071/Select_123/n2 , 
        \useone/select_1071/Select_124/n2 , \useone/select_1071/Select_125/n2 , 
        \useone/select_1071/Select_126/n2 , \useone/select_1071/Select_127/n2 , 
        \useone/n39171 , \useone/select_1071/Select_129/n2 , \useone/select_1071/Select_130/n2 , 
        \useone/select_1071/Select_131/n2 , \useone/n39167 , \useone/select_1071/Select_133/n2 , 
        \useone/select_1071/Select_134/n2 , \useone/select_1071/Select_135/n2 , 
        \useone/select_1071/Select_136/n2 , \useone/select_1071/Select_137/n2 , 
        \useone/select_1071/Select_138/n2 , \useone/select_1071/Select_139/n2 , 
        \useone/select_1071/Select_140/n2 , \useone/select_1071/Select_141/n2 , 
        \useone/select_1071/Select_142/n2 , \useone/select_1071/Select_143/n2 , 
        \useone/select_1071/Select_144/n2 , \useone/select_1071/Select_145/n2 , 
        \useone/select_1071/Select_146/n2 , \useone/select_1071/Select_147/n2 , 
        \useone/select_1071/Select_148/n2 , \useone/select_1071/Select_149/n2 , 
        \useone/select_1071/Select_150/n2 , \useone/select_1071/Select_151/n2 , 
        \useone/select_1071/Select_152/n2 , \useone/select_1071/Select_153/n2 , 
        \useone/select_1071/Select_154/n2 , \useone/select_1071/Select_155/n2 , 
        \useone/select_1071/Select_156/n2 , \useone/select_1071/Select_157/n2 , 
        \useone/select_1071/Select_158/n2 , \useone/select_1071/Select_159/n2 , 
        \useone/select_1071/Select_160/n2 , \useone/select_1071/Select_161/n2 , 
        \useone/select_1071/Select_162/n2 , \useone/select_1071/Select_163/n2 , 
        \useone/select_1071/Select_164/n2 , \useone/select_1071/Select_165/n2 , 
        \useone/select_1071/Select_166/n2 , \useone/select_1071/Select_167/n2 , 
        \useone/select_1071/Select_168/n2 , \useone/select_1071/Select_169/n2 , 
        \useone/select_1071/Select_170/n2 , \useone/select_1071/Select_171/n2 , 
        \useone/select_1071/Select_172/n2 , \useone/select_1071/Select_173/n2 , 
        \useone/select_1071/Select_174/n2 , \useone/select_1071/Select_175/n2 , 
        \useone/select_1071/Select_176/n2 , \useone/select_1071/Select_177/n2 , 
        \useone/select_1071/Select_178/n2 , \useone/select_1071/Select_179/n2 , 
        \useone/select_1071/Select_180/n2 , \useone/select_1071/Select_181/n2 , 
        \useone/select_1071/Select_182/n2 , \useone/select_1071/Select_183/n2 , 
        \useone/select_1071/Select_184/n2 , \useone/select_1071/Select_185/n2 , 
        \useone/select_1071/Select_186/n2 , \useone/select_1071/Select_187/n2 , 
        \useone/select_1071/Select_188/n2 , \useone/select_1071/Select_189/n2 , 
        \useone/select_1071/Select_190/n2 , \useone/select_1071/Select_191/n2 , 
        \useone/select_1071/Select_192/n6 , \useone/select_1071/Select_193/n2 , 
        \useone/select_1071/Select_194/n2 , \useone/select_1071/Select_195/n2 , 
        \useone/select_1071/Select_196/n2 , \useone/select_1071/Select_197/n2 , 
        \useone/select_1071/Select_198/n2 , \useone/select_1071/Select_199/n2 , 
        \useone/select_1071/Select_200/n2 , \useone/select_1071/Select_201/n2 , 
        \useone/select_1071/Select_202/n2 , \useone/select_1071/Select_203/n2 , 
        \useone/select_1071/Select_204/n2 , \useone/select_1071/Select_205/n6 , 
        \useone/select_1071/Select_206/n2 , \useone/select_1071/Select_207/n2 , 
        \useone/select_1071/Select_208/n2 , \useone/select_1071/Select_209/n2 , 
        \useone/select_1071/Select_210/n2 , \useone/select_1071/Select_211/n2 , 
        \useone/select_1071/Select_212/n2 , \useone/select_1071/Select_213/n2 , 
        \useone/select_1071/Select_214/n2 , \useone/select_1071/Select_215/n2 , 
        \useone/select_1071/Select_216/n2 , \useone/select_1071/Select_217/n2 , 
        \useone/select_1071/Select_218/n2 , \useone/select_1071/Select_219/n2 , 
        \useone/select_1071/Select_220/n2 , \useone/select_1071/Select_221/n2 , 
        \useone/select_1071/Select_222/n2 , \useone/select_1071/Select_223/n2 , 
        \useone/select_1071/Select_224/n2 , \useone/select_1071/Select_225/n2 , 
        \useone/select_1071/Select_226/n2 , \useone/select_1071/Select_227/n2 , 
        \useone/select_1071/Select_228/n2 , \useone/select_1071/Select_229/n2 , 
        \useone/select_1071/Select_230/n2 , \useone/select_1071/Select_231/n2 , 
        \useone/select_1071/Select_232/n2 , \useone/select_1071/Select_233/n2 , 
        \useone/select_1071/Select_234/n2 , \useone/select_1071/Select_235/n2 , 
        \useone/select_1071/Select_236/n2 , \useone/select_1071/Select_237/n2 , 
        \useone/select_1071/Select_238/n2 , \useone/select_1071/Select_239/n2 , 
        \useone/select_1071/Select_240/n2 , \useone/select_1071/Select_241/n2 , 
        \useone/select_1071/Select_242/n2 , \useone/select_1071/Select_243/n2 , 
        \useone/select_1071/Select_244/n2 , \useone/select_1071/Select_245/n2 , 
        \useone/select_1071/Select_246/n2 , \useone/select_1071/Select_247/n2 , 
        \useone/select_1071/Select_248/n2 , \useone/select_1071/Select_249/n2 , 
        \useone/select_1071/Select_250/n2 , \useone/select_1071/Select_251/n2 , 
        \useone/select_1071/Select_252/n2 , \useone/select_1071/Select_253/n2 , 
        \useone/select_1071/Select_254/n2 , \useone/select_1071/Select_255/n2 , 
        \useuart/n844 , \useuart/r_SM_Main[2] , \useuart/n634 , \useuart/n848 , 
        ceg_net79, \useuart/r_SM_Main[1] , ceg_net77, \useuart/n960 , 
        \useuart/n840 , \useuart/n708 , \useuart/n711 , \useuart/n714 , 
        \useuart/n717 , \useuart/n720 , \useuart/n723 , \useuart/n726 , 
        \useuart/n729 , \useuart/n732 , \useuart/n735 , \useuart/n738 , 
        \useuart/n741 , \useuart/n802 , \useuart/n806 , \data_chunk[1] , 
        \data_chunk[2] , \data_chunk[3] , \data_chunk[4] , \data_chunk[5] , 
        \data_chunk[6] , \data_chunk[7] , \useuart/n836 , \useuart/LessThan_9/n26 , 
        \useuart/n942 , n827, n826, n825, n824, n823, n822, n821, 
        n3421, n3422, n3424, n3425, n3427, n3428, n3430, n3431, 
        n3433, n3434, n3436, n3437, n3439, n3440, n3442, n3443, 
        n3445, n3446, n3448, n3449, n3451, n3452, n3454, n3455, 
        n3457, n3458, n3460, n3461, n3463, n3464, n3466, n3467, 
        n3469, n3470, n3472, n3473, n3475, n3476, n3478, n3479, 
        n3481, n3482, n3484, n3485, n3487, n3488, n3490, n3491, 
        n3493, n3494, n3496, n3497, n3499, n3500, n3502, n3503, 
        n3505, n3506, n3508, n3509, n3511, n3512, n3515, n3518, 
        n3521, n3524, n3527, n3530, n3533, n3536, n3539, n3542, 
        n3545, n3548, n3551, n3554, n3557, n3560, n3563, n3566, 
        n3569, n3572, n3575, n3578, n3581, n3584, n3587, n3590, 
        n3593, n3596, n3599, n3602, n3605, n3608, n3611, n3614, 
        n3617, n3620, n3623, n3626, n3629, n3632, n3635, n3638, 
        n3641, n3644, n3647, n3650, n3653, n3656, n3659, n3662, 
        n3665, n3668, n3671, n3674, n3677, n3680, n3683, n3686, 
        n3689, n3692, n3695, n3698, n3701, n3704, n3707, n3710, 
        n3713, n3716, n3719, n3722, n3725, n3728, n3731, n3734, 
        n3737, n3740, n3743, n3746, n3749, n3752, n3755, n3758, 
        n3761, n3764, n3767, n3770, n3773, n3776, n3779, n3782, 
        n3785, n3788, n3791, n3793, n3795, n3797, n3799, n3801, 
        n3803, n3805, n3807, n3809, n3811, n3813, n3815, n3817, 
        n3819, n3821, n3823, n3825, n3827, n3829, n3831, n3833, 
        n3835, n3837, n3839, n3841, n3843, n3845, n3847, n3849, 
        n3851, n3853, \clk~O , \useone/equal_1067/n7 , n3857, n3858, 
        n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, 
        n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, 
        n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, 
        n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, 
        n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, 
        n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, 
        n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, 
        n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, 
        n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, 
        n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, 
        n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, 
        n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, 
        n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, 
        n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, 
        n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, 
        n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, 
        n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, 
        n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, 
        n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, 
        n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, 
        n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, 
        n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, 
        n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
        n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, 
        n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, 
        n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, 
        n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, 
        n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, 
        n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, 
        n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
        n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, 
        n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, 
        n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, 
        n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, 
        n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, 
        n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, 
        n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, 
        n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, 
        n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, 
        n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
        n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, 
        n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, 
        n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, 
        n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, 
        n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
        n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, 
        n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, 
        n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, 
        n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, 
        n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, 
        n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, 
        n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, 
        n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, 
        n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, 
        n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, 
        n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, 
        n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, 
        n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, 
        n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, 
        n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, 
        n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, 
        n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, 
        n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
        n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, 
        n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, 
        n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, 
        n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, 
        n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, 
        n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, 
        n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, 
        n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, 
        n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, 
        n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
        n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, 
        n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, 
        n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, 
        n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, 
        n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, 
        n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, 
        n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, 
        n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, 
        n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, 
        n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, 
        n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, 
        n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, 
        n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, 
        n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, 
        n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, 
        n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, 
        n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, 
        n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, 
        n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, 
        n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, 
        n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, 
        n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, 
        n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, 
        n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, 
        n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, 
        n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, 
        n4651, n4652, n4653;
    
    EFX_FF \chunk_index[0]~FF  (.D(\chunk_index[0] ), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\chunk_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \chunk_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \chunk_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \chunk_index[0]~FF .SR_POLARITY = 1'b1;
    defparam \chunk_index[0]~FF .D_POLARITY = 1'b0;
    defparam \chunk_index[0]~FF .SR_SYNC = 1'b0;
    defparam \chunk_index[0]~FF .SR_VALUE = 1'b0;
    defparam \chunk_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \done~FF  (.D(1'b1), .CE(ceg_net85), .CLK(\clk~O ), .SR(rst), 
           .Q(done)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \done~FF .CLK_POLARITY = 1'b1;
    defparam \done~FF .CE_POLARITY = 1'b1;
    defparam \done~FF .SR_POLARITY = 1'b1;
    defparam \done~FF .D_POLARITY = 1'b1;
    defparam \done~FF .SR_SYNC = 1'b0;
    defparam \done~FF .SR_VALUE = 1'b0;
    defparam \done~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \tx_valid~FF  (.D(\state[1] ), .CE(ceg_net86), .CLK(\clk~O ), 
           .SR(rst), .Q(tx_valid)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \tx_valid~FF .CLK_POLARITY = 1'b1;
    defparam \tx_valid~FF .CE_POLARITY = 1'b0;
    defparam \tx_valid~FF .SR_POLARITY = 1'b1;
    defparam \tx_valid~FF .D_POLARITY = 1'b0;
    defparam \tx_valid~FF .SR_SYNC = 1'b0;
    defparam \tx_valid~FF .SR_VALUE = 1'b0;
    defparam \tx_valid~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \state[0]~FF  (.D(n869_2), .CE(ceg_net99), .CLK(\clk~O ), .SR(rst), 
           .Q(\state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \state[0]~FF .CE_POLARITY = 1'b0;
    defparam \state[0]~FF .SR_POLARITY = 1'b1;
    defparam \state[0]~FF .D_POLARITY = 1'b1;
    defparam \state[0]~FF .SR_SYNC = 1'b0;
    defparam \state[0]~FF .SR_VALUE = 1'b0;
    defparam \state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_chunk[0]~FF  (.D(n828_2), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\data_chunk[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \data_chunk[0]~FF .CLK_POLARITY = 1'b1;
    defparam \data_chunk[0]~FF .CE_POLARITY = 1'b0;
    defparam \data_chunk[0]~FF .SR_POLARITY = 1'b1;
    defparam \data_chunk[0]~FF .D_POLARITY = 1'b1;
    defparam \data_chunk[0]~FF .SR_SYNC = 1'b0;
    defparam \data_chunk[0]~FF .SR_VALUE = 1'b0;
    defparam \data_chunk[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/state[0]~FF  (.D(\useone/select_1072/Select_0/n5 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/state[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/state[0]~FF .D_POLARITY = 1'b1;
    defparam \useone/state[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/state[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[0]~FF  (.D(n22), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[0]~FF  (.D(\useone/a[0] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[0]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[0]~FF  (.D(\useone/b[0] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[0]~FF  (.D(\useone/c[0] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[0]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[0]~FF  (.D(n20), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[0]~FF  (.D(\useone/e[0] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[0]~FF  (.D(\useone/f[0] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[0]~FF  (.D(\useone/g[0] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[0]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/round_flag[0]~FF  (.D(\useone/round_flag[0] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/round_flag[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/round_flag[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/round_flag[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/round_flag[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/round_flag[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/round_flag[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/round_flag[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/round_flag[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[0]~FF  (.D(n24), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[0]~FF  (.D(n26), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[0]~FF  (.D(n28), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[0]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[0]~FF  (.D(n30), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[0]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[0]~FF  (.D(n32), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[0]~FF  (.D(n34), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[0]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[0]~FF  (.D(n36), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[0]~FF  (.D(n38), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[0]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[0]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[0]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[0]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[0]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \hashdone~FF  (.D(1'b1), .CE(\useone/equal_1069/n7 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(hashdone)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \hashdone~FF .CLK_POLARITY = 1'b1;
    defparam \hashdone~FF .CE_POLARITY = 1'b0;
    defparam \hashdone~FF .SR_POLARITY = 1'b1;
    defparam \hashdone~FF .D_POLARITY = 1'b1;
    defparam \hashdone~FF .SR_SYNC = 1'b1;
    defparam \hashdone~FF .SR_VALUE = 1'b0;
    defparam \hashdone~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[0]~FF  (.D(\useone/select_1071/Select_0/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[0]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[0]~FF .CE_POLARITY = 1'b1;
    defparam \signature[0]~FF .SR_POLARITY = 1'b1;
    defparam \signature[0]~FF .D_POLARITY = 1'b1;
    defparam \signature[0]~FF .SR_SYNC = 1'b1;
    defparam \signature[0]~FF .SR_VALUE = 1'b0;
    defparam \signature[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/state[1]~FF  (.D(\useone/select_1072/Select_1/n8 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/state[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/state[1]~FF .D_POLARITY = 1'b1;
    defparam \useone/state[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/state[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/state[2]~FF  (.D(\useone/n39302 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/state[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/state[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/state[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/state[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/state[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[1]~FF  (.D(n1408), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[2]~FF  (.D(n1406), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[2]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[3]~FF  (.D(n1404), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[4]~FF  (.D(n1402), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[5]~FF  (.D(n1400), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[6]~FF  (.D(n1398), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[7]~FF  (.D(n1396), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[8]~FF  (.D(n1394), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[9]~FF  (.D(n1392), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[9]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[10]~FF  (.D(n1390), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[10]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[11]~FF  (.D(n1388), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[12]~FF  (.D(n1386), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[12]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[13]~FF  (.D(n1384), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[13]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[14]~FF  (.D(n1382), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[15]~FF  (.D(n1380), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[15]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[16]~FF  (.D(n1378), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[17]~FF  (.D(n1376), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[17]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[18]~FF  (.D(n1374), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[18]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[19]~FF  (.D(n1372), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[20]~FF  (.D(n1370), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[21]~FF  (.D(n1368), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[22]~FF  (.D(n1366), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[23]~FF  (.D(n1364), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[24]~FF  (.D(n1362), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[24]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[25]~FF  (.D(n1360), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[25]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[26]~FF  (.D(n1358), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[27]~FF  (.D(n1356), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[28]~FF  (.D(n1354), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[28]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[29]~FF  (.D(n1352), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[29]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[30]~FF  (.D(n1350), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[30]~FF .D_POLARITY = 1'b0;
    defparam \useone/a[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/a[31]~FF  (.D(n1349), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/a[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/a[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/a[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/a[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/a[31]~FF .D_POLARITY = 1'b1;
    defparam \useone/a[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/a[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/a[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[1]~FF  (.D(\useone/a[1] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[2]~FF  (.D(\useone/a[2] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[3]~FF  (.D(\useone/a[3] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[4]~FF  (.D(\useone/a[4] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[5]~FF  (.D(\useone/a[5] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[6]~FF  (.D(\useone/a[6] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[7]~FF  (.D(\useone/a[7] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[7]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[8]~FF  (.D(\useone/a[8] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[9]~FF  (.D(\useone/a[9] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/b[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[9]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[10]~FF  (.D(\useone/a[10] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[10]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[11]~FF  (.D(\useone/a[11] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[11]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[12]~FF  (.D(\useone/a[12] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[12]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[13]~FF  (.D(\useone/a[13] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[13]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[14]~FF  (.D(\useone/a[14] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[15]~FF  (.D(\useone/a[15] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[15]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[16]~FF  (.D(\useone/a[16] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[16]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[17]~FF  (.D(\useone/a[17] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[18]~FF  (.D(\useone/a[18] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[18]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[19]~FF  (.D(\useone/a[19] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[20]~FF  (.D(\useone/a[20] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[21]~FF  (.D(\useone/a[21] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[21]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[22]~FF  (.D(\useone/a[22] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[22]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[23]~FF  (.D(\useone/a[23] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[24]~FF  (.D(\useone/a[24] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[25]~FF  (.D(\useone/a[25] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[25]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[26]~FF  (.D(\useone/a[26] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[27]~FF  (.D(\useone/a[27] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[27]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[28]~FF  (.D(\useone/a[28] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[29]~FF  (.D(\useone/a[29] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/b[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[30]~FF  (.D(\useone/a[30] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[30]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/b[31]~FF  (.D(\useone/a[31] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/b[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/b[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/b[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/b[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/b[31]~FF .D_POLARITY = 1'b0;
    defparam \useone/b[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/b[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/b[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[1]~FF  (.D(\useone/b[1] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[2]~FF  (.D(\useone/b[2] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[2]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[3]~FF  (.D(\useone/b[3] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[4]~FF  (.D(\useone/b[4] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[4]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[5]~FF  (.D(\useone/b[5] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[6]~FF  (.D(\useone/b[6] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[7]~FF  (.D(\useone/b[7] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[7]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[8]~FF  (.D(\useone/b[8] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[8]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[9]~FF  (.D(\useone/b[9] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/c[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[9]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[10]~FF  (.D(\useone/b[10] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[10]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[11]~FF  (.D(\useone/b[11] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[11]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[12]~FF  (.D(\useone/b[12] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[13]~FF  (.D(\useone/b[13] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[13]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[14]~FF  (.D(\useone/b[14] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[15]~FF  (.D(\useone/b[15] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[15]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[16]~FF  (.D(\useone/b[16] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[17]~FF  (.D(\useone/b[17] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[17]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[18]~FF  (.D(\useone/b[18] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[18]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[19]~FF  (.D(\useone/b[19] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[20]~FF  (.D(\useone/b[20] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[21]~FF  (.D(\useone/b[21] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[22]~FF  (.D(\useone/b[22] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[23]~FF  (.D(\useone/b[23] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[24]~FF  (.D(\useone/b[24] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[25]~FF  (.D(\useone/b[25] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[25]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[26]~FF  (.D(\useone/b[26] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[26]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[27]~FF  (.D(\useone/b[27] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[27]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[28]~FF  (.D(\useone/b[28] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[28]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[29]~FF  (.D(\useone/b[29] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[30]~FF  (.D(\useone/b[30] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[30]~FF .D_POLARITY = 1'b1;
    defparam \useone/c[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/c[31]~FF  (.D(\useone/b[31] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/c[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/c[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/c[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/c[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/c[31]~FF .D_POLARITY = 1'b0;
    defparam \useone/c[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/c[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/c[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[1]~FF  (.D(\useone/c[1] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[1]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[2]~FF  (.D(\useone/c[2] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[3]~FF  (.D(\useone/c[3] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[3]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[4]~FF  (.D(\useone/c[4] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[5]~FF  (.D(\useone/c[5] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[5]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[6]~FF  (.D(\useone/c[6] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[7]~FF  (.D(\useone/c[7] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[8]~FF  (.D(\useone/c[8] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[9]~FF  (.D(\useone/c[9] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/d[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[9]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[10]~FF  (.D(\useone/c[10] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[10]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[11]~FF  (.D(\useone/c[11] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[12]~FF  (.D(\useone/c[12] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[12]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[13]~FF  (.D(\useone/c[13] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[13]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[14]~FF  (.D(\useone/c[14] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[14]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[15]~FF  (.D(\useone/c[15] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[15]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[16]~FF  (.D(\useone/c[16] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[17]~FF  (.D(\useone/c[17] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[17]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[18]~FF  (.D(\useone/c[18] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[18]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[19]~FF  (.D(\useone/c[19] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[19]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[20]~FF  (.D(\useone/c[20] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[21]~FF  (.D(\useone/c[21] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[21]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[22]~FF  (.D(\useone/c[22] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[23]~FF  (.D(\useone/c[23] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[24]~FF  (.D(\useone/c[24] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[25]~FF  (.D(\useone/c[25] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[25]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[26]~FF  (.D(\useone/c[26] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[27]~FF  (.D(\useone/c[27] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[28]~FF  (.D(\useone/c[28] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[29]~FF  (.D(\useone/c[29] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[30]~FF  (.D(\useone/c[30] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[30]~FF .D_POLARITY = 1'b1;
    defparam \useone/d[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/d[31]~FF  (.D(\useone/c[31] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/d[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/d[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/d[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/d[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/d[31]~FF .D_POLARITY = 1'b0;
    defparam \useone/d[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/d[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/d[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[1]~FF  (.D(n1469), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[2]~FF  (.D(n1467), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[2]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[3]~FF  (.D(n1465), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[3]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[4]~FF  (.D(n1463), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[4]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[5]~FF  (.D(n1461), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[6]~FF  (.D(n1459), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[7]~FF  (.D(n1457), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[8]~FF  (.D(n1455), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[9]~FF  (.D(n1453), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[9]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[10]~FF  (.D(n1451), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[10]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[11]~FF  (.D(n1449), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[12]~FF  (.D(n1447), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[13]~FF  (.D(n1445), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[13]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[14]~FF  (.D(n1443), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[15]~FF  (.D(n1441), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[15]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[16]~FF  (.D(n1439), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[16]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[17]~FF  (.D(n1437), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[18]~FF  (.D(n1435), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[18]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[19]~FF  (.D(n1433), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[20]~FF  (.D(n1431), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[21]~FF  (.D(n1429), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[22]~FF  (.D(n1427), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[23]~FF  (.D(n1425), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[24]~FF  (.D(n1423), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[25]~FF  (.D(n1421), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[25]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[26]~FF  (.D(n1419), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[27]~FF  (.D(n1417), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[27]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[28]~FF  (.D(n1415), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[29]~FF  (.D(n1413), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[30]~FF  (.D(n1411), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[30]~FF .D_POLARITY = 1'b0;
    defparam \useone/e[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/e[31]~FF  (.D(n1410), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/e[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/e[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/e[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/e[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/e[31]~FF .D_POLARITY = 1'b1;
    defparam \useone/e[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/e[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/e[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[1]~FF  (.D(\useone/e[1] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[2]~FF  (.D(\useone/e[2] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[3]~FF  (.D(\useone/e[3] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[4]~FF  (.D(\useone/e[4] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[4]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[5]~FF  (.D(\useone/e[5] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[6]~FF  (.D(\useone/e[6] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[7]~FF  (.D(\useone/e[7] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[7]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[8]~FF  (.D(\useone/e[8] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[9]~FF  (.D(\useone/e[9] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/f[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[9]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[10]~FF  (.D(\useone/e[10] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[10]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[11]~FF  (.D(\useone/e[11] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[11]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[12]~FF  (.D(\useone/e[12] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[13]~FF  (.D(\useone/e[13] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[13]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[14]~FF  (.D(\useone/e[14] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[14]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[15]~FF  (.D(\useone/e[15] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[15]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[16]~FF  (.D(\useone/e[16] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[17]~FF  (.D(\useone/e[17] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[18]~FF  (.D(\useone/e[18] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[18]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[19]~FF  (.D(\useone/e[19] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[20]~FF  (.D(\useone/e[20] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[21]~FF  (.D(\useone/e[21] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[22]~FF  (.D(\useone/e[22] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[23]~FF  (.D(\useone/e[23] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[24]~FF  (.D(\useone/e[24] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[24]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[25]~FF  (.D(\useone/e[25] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[25]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[26]~FF  (.D(\useone/e[26] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[27]~FF  (.D(\useone/e[27] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[28]~FF  (.D(\useone/e[28] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[28]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[29]~FF  (.D(\useone/e[29] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/f[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[30]~FF  (.D(\useone/e[30] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[30]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/f[31]~FF  (.D(\useone/e[31] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/f[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/f[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/f[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/f[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/f[31]~FF .D_POLARITY = 1'b0;
    defparam \useone/f[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/f[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/f[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[1]~FF  (.D(\useone/f[1] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[2]~FF  (.D(\useone/f[2] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[2]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[3]~FF  (.D(\useone/f[3] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[4]~FF  (.D(\useone/f[4] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[5]~FF  (.D(\useone/f[5] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[6]~FF  (.D(\useone/f[6] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[6]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[7]~FF  (.D(\useone/f[7] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[8]~FF  (.D(\useone/f[8] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[8]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[9]~FF  (.D(\useone/f[9] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/g[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[9]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[10]~FF  (.D(\useone/f[10] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[10]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[11]~FF  (.D(\useone/f[11] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[12]~FF  (.D(\useone/f[12] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[13]~FF  (.D(\useone/f[13] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[13]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[14]~FF  (.D(\useone/f[14] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[14]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[15]~FF  (.D(\useone/f[15] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[15]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[16]~FF  (.D(\useone/f[16] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[16]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[17]~FF  (.D(\useone/f[17] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[18]~FF  (.D(\useone/f[18] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[18]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[19]~FF  (.D(\useone/f[19] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[19]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[20]~FF  (.D(\useone/f[20] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[21]~FF  (.D(\useone/f[21] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[22]~FF  (.D(\useone/f[22] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[23]~FF  (.D(\useone/f[23] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[23]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[24]~FF  (.D(\useone/f[24] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[24]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[25]~FF  (.D(\useone/f[25] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[25]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[26]~FF  (.D(\useone/f[26] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[26]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[27]~FF  (.D(\useone/f[27] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[27]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[28]~FF  (.D(\useone/f[28] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[28]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[29]~FF  (.D(\useone/f[29] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[30]~FF  (.D(\useone/f[30] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[30]~FF .D_POLARITY = 1'b1;
    defparam \useone/g[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/g[31]~FF  (.D(\useone/f[31] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/g[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/g[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/g[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/g[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/g[31]~FF .D_POLARITY = 1'b0;
    defparam \useone/g[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/g[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/g[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[1]~FF  (.D(\useone/g[1] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[2]~FF  (.D(\useone/g[2] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[3]~FF  (.D(\useone/g[3] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[4]~FF  (.D(\useone/g[4] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[4]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[5]~FF  (.D(\useone/g[5] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[6]~FF  (.D(\useone/g[6] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[6]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[7]~FF  (.D(\useone/g[7] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[7]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[8]~FF  (.D(\useone/g[8] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[9]~FF  (.D(\useone/g[9] ), .CE(\useone/n144202 ), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\useone/h[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[9]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[10]~FF  (.D(\useone/g[10] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[10]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[11]~FF  (.D(\useone/g[11] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[12]~FF  (.D(\useone/g[12] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[13]~FF  (.D(\useone/g[13] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[13]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[14]~FF  (.D(\useone/g[14] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[14]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[15]~FF  (.D(\useone/g[15] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[15]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[16]~FF  (.D(\useone/g[16] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[17]~FF  (.D(\useone/g[17] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[18]~FF  (.D(\useone/g[18] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[18]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[19]~FF  (.D(\useone/g[19] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[19]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[20]~FF  (.D(\useone/g[20] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[21]~FF  (.D(\useone/g[21] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[21]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[22]~FF  (.D(\useone/g[22] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[22]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[23]~FF  (.D(\useone/g[23] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[24]~FF  (.D(\useone/g[24] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[24]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[25]~FF  (.D(\useone/g[25] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[25]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[26]~FF  (.D(\useone/g[26] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[26]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[27]~FF  (.D(\useone/g[27] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[27]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[28]~FF  (.D(\useone/g[28] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[28]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[29]~FF  (.D(\useone/g[29] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[30]~FF  (.D(\useone/g[30] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[30]~FF .D_POLARITY = 1'b0;
    defparam \useone/h[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/h[31]~FF  (.D(\useone/g[31] ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/h[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/h[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/h[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/h[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/h[31]~FF .D_POLARITY = 1'b1;
    defparam \useone/h[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/h[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/h[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/round_flag[1]~FF  (.D(\useone/n46233 ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/round_flag[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/round_flag[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/round_flag[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/round_flag[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/round_flag[1]~FF .D_POLARITY = 1'b1;
    defparam \useone/round_flag[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/round_flag[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/round_flag[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/round_flag[2]~FF  (.D(\useone/n46238 ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/round_flag[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/round_flag[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/round_flag[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/round_flag[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/round_flag[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/round_flag[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/round_flag[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/round_flag[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/round_flag[3]~FF  (.D(\useone/n46243 ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/round_flag[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/round_flag[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/round_flag[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/round_flag[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/round_flag[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/round_flag[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/round_flag[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/round_flag[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/round_flag[4]~FF  (.D(\useone/n46248 ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/round_flag[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/round_flag[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/round_flag[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/round_flag[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/round_flag[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/round_flag[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/round_flag[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/round_flag[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/round_flag[5]~FF  (.D(\useone/n46253 ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/round_flag[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/round_flag[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/round_flag[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/round_flag[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/round_flag[5]~FF .D_POLARITY = 1'b1;
    defparam \useone/round_flag[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/round_flag[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/round_flag[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/round_flag[6]~FF  (.D(\useone/n46258 ), .CE(\useone/n144202 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/round_flag[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/round_flag[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/round_flag[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/round_flag[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/round_flag[6]~FF .D_POLARITY = 1'b1;
    defparam \useone/round_flag[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/round_flag[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/round_flag[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[1]~FF  (.D(n1347), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[2]~FF  (.D(n1345), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[2]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[3]~FF  (.D(n1343), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[4]~FF  (.D(n1341), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[5]~FF  (.D(n1339), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[6]~FF  (.D(n1337), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[7]~FF  (.D(n1335), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[8]~FF  (.D(n1333), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[9]~FF  (.D(n1331), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[9]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[10]~FF  (.D(n1329), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[10]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[11]~FF  (.D(n1327), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[12]~FF  (.D(n1325), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[12]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[13]~FF  (.D(n1323), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[13]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[14]~FF  (.D(n1321), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[15]~FF  (.D(n1319), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[15]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[16]~FF  (.D(n1317), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[17]~FF  (.D(n1315), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[17]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[18]~FF  (.D(n1313), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[18]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[19]~FF  (.D(n1311), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[20]~FF  (.D(n1309), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[21]~FF  (.D(n1307), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[22]~FF  (.D(n1305), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[23]~FF  (.D(n1303), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[24]~FF  (.D(n1301), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[24]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[25]~FF  (.D(n1299), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[25]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[26]~FF  (.D(n1297), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[27]~FF  (.D(n1295), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[28]~FF  (.D(n1293), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[28]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[29]~FF  (.D(n1291), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[29]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[30]~FF  (.D(n1289), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[30]~FF .D_POLARITY = 1'b0;
    defparam \useone/H0[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H0[31]~FF  (.D(n1288), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H0[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H0[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H0[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H0[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H0[31]~FF .D_POLARITY = 1'b1;
    defparam \useone/H0[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/H0[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/H0[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[1]~FF  (.D(n1286), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[1]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[2]~FF  (.D(n1284), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[2]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[3]~FF  (.D(n1282), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[4]~FF  (.D(n1280), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[5]~FF  (.D(n1278), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[5]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[6]~FF  (.D(n1276), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[6]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[7]~FF  (.D(n1274), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[7]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[8]~FF  (.D(n1272), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[9]~FF  (.D(n1270), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[9]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[10]~FF  (.D(n1268), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[10]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[11]~FF  (.D(n1266), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[11]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[12]~FF  (.D(n1264), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[12]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[13]~FF  (.D(n1262), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[13]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[14]~FF  (.D(n1260), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[14]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[15]~FF  (.D(n1258), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[15]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[16]~FF  (.D(n1256), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[17]~FF  (.D(n1254), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[18]~FF  (.D(n1252), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[18]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[19]~FF  (.D(n1250), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[19]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[20]~FF  (.D(n1248), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[21]~FF  (.D(n1246), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[21]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[22]~FF  (.D(n1244), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[22]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[23]~FF  (.D(n1242), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[24]~FF  (.D(n1240), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[25]~FF  (.D(n1238), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[25]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[26]~FF  (.D(n1236), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[27]~FF  (.D(n1234), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[28]~FF  (.D(n1232), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[29]~FF  (.D(n1230), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[29]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[30]~FF  (.D(n1228), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[30]~FF .D_POLARITY = 1'b1;
    defparam \useone/H1[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H1[31]~FF  (.D(n1227), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H1[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H1[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H1[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H1[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H1[31]~FF .D_POLARITY = 1'b0;
    defparam \useone/H1[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/H1[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/H1[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[1]~FF  (.D(n1225), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[2]~FF  (.D(n1223), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[3]~FF  (.D(n1221), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[3]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[4]~FF  (.D(n1219), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[4]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[5]~FF  (.D(n1217), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[6]~FF  (.D(n1215), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[7]~FF  (.D(n1213), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[8]~FF  (.D(n1211), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[8]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[9]~FF  (.D(n1209), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[9]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[10]~FF  (.D(n1207), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[10]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[11]~FF  (.D(n1205), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[12]~FF  (.D(n1203), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[13]~FF  (.D(n1201), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[13]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[14]~FF  (.D(n1199), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[15]~FF  (.D(n1197), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[15]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[16]~FF  (.D(n1195), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[16]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[17]~FF  (.D(n1193), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[18]~FF  (.D(n1191), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[18]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[19]~FF  (.D(n1189), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[20]~FF  (.D(n1187), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[21]~FF  (.D(n1185), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[21]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[22]~FF  (.D(n1183), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[22]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[23]~FF  (.D(n1181), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[24]~FF  (.D(n1179), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[24]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[25]~FF  (.D(n1177), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[25]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[26]~FF  (.D(n1175), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[26]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[27]~FF  (.D(n1173), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[28]~FF  (.D(n1171), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[29]~FF  (.D(n1169), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[29]~FF .D_POLARITY = 1'b0;
    defparam \useone/H2[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[30]~FF  (.D(n1167), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[30]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H2[31]~FF  (.D(n1166), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H2[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H2[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H2[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H2[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H2[31]~FF .D_POLARITY = 1'b1;
    defparam \useone/H2[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/H2[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/H2[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[1]~FF  (.D(n1164), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[2]~FF  (.D(n1162), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[3]~FF  (.D(n1160), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[3]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[4]~FF  (.D(n1158), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[4]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[5]~FF  (.D(n1156), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[6]~FF  (.D(n1154), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[6]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[7]~FF  (.D(n1152), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[8]~FF  (.D(n1150), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[8]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[9]~FF  (.D(n1148), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[9]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[10]~FF  (.D(n1146), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[10]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[11]~FF  (.D(n1144), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[12]~FF  (.D(n1142), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[13]~FF  (.D(n1140), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[13]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[14]~FF  (.D(n1138), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[15]~FF  (.D(n1136), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[15]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[16]~FF  (.D(n1134), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[17]~FF  (.D(n1132), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[18]~FF  (.D(n1130), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[18]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[19]~FF  (.D(n1128), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[20]~FF  (.D(n1126), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[21]~FF  (.D(n1124), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[22]~FF  (.D(n1122), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[22]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[23]~FF  (.D(n1120), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[24]~FF  (.D(n1118), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[25]~FF  (.D(n1116), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[25]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[26]~FF  (.D(n1114), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[26]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[27]~FF  (.D(n1112), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[27]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[28]~FF  (.D(n1110), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[28]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[29]~FF  (.D(n1108), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[29]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[30]~FF  (.D(n1106), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[30]~FF .D_POLARITY = 1'b1;
    defparam \useone/H3[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H3[31]~FF  (.D(n1105), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H3[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H3[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H3[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H3[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H3[31]~FF .D_POLARITY = 1'b0;
    defparam \useone/H3[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/H3[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/H3[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[1]~FF  (.D(n1103), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[2]~FF  (.D(n1101), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[2]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[3]~FF  (.D(n1099), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[3]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[4]~FF  (.D(n1097), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[4]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[5]~FF  (.D(n1095), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[6]~FF  (.D(n1093), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[6]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[7]~FF  (.D(n1091), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[8]~FF  (.D(n1089), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[9]~FF  (.D(n1087), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[9]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[10]~FF  (.D(n1085), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[10]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[11]~FF  (.D(n1083), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[11]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[12]~FF  (.D(n1081), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[13]~FF  (.D(n1079), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[13]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[14]~FF  (.D(n1077), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[15]~FF  (.D(n1075), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[15]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[16]~FF  (.D(n1073), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[16]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[17]~FF  (.D(n1071), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[18]~FF  (.D(n1069), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[18]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[19]~FF  (.D(n1067), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[19]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[20]~FF  (.D(n1065), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[21]~FF  (.D(n1063), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[22]~FF  (.D(n1061), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[23]~FF  (.D(n1059), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[24]~FF  (.D(n1057), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[25]~FF  (.D(n1055), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[25]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[26]~FF  (.D(n1053), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[27]~FF  (.D(n1051), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[27]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[28]~FF  (.D(n1049), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[29]~FF  (.D(n1047), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[30]~FF  (.D(n1045), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[30]~FF .D_POLARITY = 1'b0;
    defparam \useone/H4[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H4[31]~FF  (.D(n1044), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H4[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H4[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H4[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H4[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H4[31]~FF .D_POLARITY = 1'b1;
    defparam \useone/H4[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/H4[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/H4[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[1]~FF  (.D(n1042), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[1]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[2]~FF  (.D(n1040), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[2]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[3]~FF  (.D(n1038), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[3]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[4]~FF  (.D(n1036), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[5]~FF  (.D(n1034), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[5]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[6]~FF  (.D(n1032), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[6]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[7]~FF  (.D(n1030), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[7]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[8]~FF  (.D(n1028), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[8]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[9]~FF  (.D(n1026), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[9]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[10]~FF  (.D(n1024), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[10]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[11]~FF  (.D(n1022), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[11]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[12]~FF  (.D(n1020), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[12]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[13]~FF  (.D(n1018), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[13]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[14]~FF  (.D(n1016), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[15]~FF  (.D(n1014), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[15]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[16]~FF  (.D(n1012), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[17]~FF  (.D(n1010), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[17]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[18]~FF  (.D(n1008), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[18]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[19]~FF  (.D(n1006), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[19]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[20]~FF  (.D(n1004), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[21]~FF  (.D(n1002), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[22]~FF  (.D(n1000), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[23]~FF  (.D(n998), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[23]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[24]~FF  (.D(n996), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[25]~FF  (.D(n994), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[25]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[26]~FF  (.D(n992), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[27]~FF  (.D(n990), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[28]~FF  (.D(n988), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[29]~FF  (.D(n986), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[30]~FF  (.D(n984), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[30]~FF .D_POLARITY = 1'b1;
    defparam \useone/H5[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H5[31]~FF  (.D(n983), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H5[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H5[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H5[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H5[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H5[31]~FF .D_POLARITY = 1'b0;
    defparam \useone/H5[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/H5[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/H5[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[1]~FF  (.D(n981), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[1]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[2]~FF  (.D(n979), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[3]~FF  (.D(n977), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[3]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[4]~FF  (.D(n975), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[4]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[5]~FF  (.D(n973), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[5]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[6]~FF  (.D(n971), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[6]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[7]~FF  (.D(n969), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[7]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[8]~FF  (.D(n967), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[8]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[9]~FF  (.D(n965), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[9]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[10]~FF  (.D(n963), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[10]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[11]~FF  (.D(n961), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[11]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[12]~FF  (.D(n959), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[12]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[13]~FF  (.D(n957), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[13]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[14]~FF  (.D(n955), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[15]~FF  (.D(n953), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[15]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[16]~FF  (.D(n951), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[16]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[17]~FF  (.D(n949), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[17]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[18]~FF  (.D(n947), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[18]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[19]~FF  (.D(n945), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[19]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[20]~FF  (.D(n943), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[21]~FF  (.D(n941), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[21]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[22]~FF  (.D(n939), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[22]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[23]~FF  (.D(n937), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[23]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[24]~FF  (.D(n935), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[25]~FF  (.D(n933), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[25]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[26]~FF  (.D(n931), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[26]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[27]~FF  (.D(n929), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[28]~FF  (.D(n927), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/H6[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[29]~FF  (.D(n925), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[30]~FF  (.D(n923), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[30]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H6[31]~FF  (.D(n922), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H6[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H6[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H6[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H6[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H6[31]~FF .D_POLARITY = 1'b1;
    defparam \useone/H6[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/H6[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/H6[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[1]~FF  (.D(n920), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[1]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[1]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[1]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[1]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[1]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[2]~FF  (.D(n918), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[2]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[2]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[2]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[2]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[2]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[3]~FF  (.D(n916), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[3]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[3]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[3]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[3]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[3]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[4]~FF  (.D(n914), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[4]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[4]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[4]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[4]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[4]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[5]~FF  (.D(n912), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[5]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[5]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[5]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[5]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[5]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[6]~FF  (.D(n910), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[6]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[6]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[6]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[6]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[6]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[7]~FF  (.D(n908), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[7]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[7]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[7]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[7]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[7]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[8]~FF  (.D(n906), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[8]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[8]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[8]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[8]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[8]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[9]~FF  (.D(n904), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[9]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[9]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[9]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[9]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[9]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[10]~FF  (.D(n902), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[10]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[10]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[10]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[10]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[10]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[11]~FF  (.D(n900), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[11]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[11]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[11]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[11]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[11]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[12]~FF  (.D(n898), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[12]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[12]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[12]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[12]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[12]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[13]~FF  (.D(n896), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[13]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[13]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[13]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[13]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[13]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[13]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[14]~FF  (.D(n894), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[14]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[14]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[14]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[14]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[14]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[14]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[15]~FF  (.D(n892), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[15]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[15]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[15]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[15]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[15]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[15]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[16]~FF  (.D(n890), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[16]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[16]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[16]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[16]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[16]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[16]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[17]~FF  (.D(n888), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[17]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[17]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[17]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[17]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[17]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[17]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[18]~FF  (.D(n886), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[18]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[18]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[18]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[18]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[18]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[18]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[19]~FF  (.D(n884), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[19]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[19]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[19]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[19]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[19]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[19]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[20]~FF  (.D(n882), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[20]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[20]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[20]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[20]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[20]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[20]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[21]~FF  (.D(n880), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[21]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[21]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[21]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[21]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[21]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[21]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[22]~FF  (.D(n878), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[22]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[22]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[22]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[22]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[22]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[22]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[23]~FF  (.D(n876), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[23]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[23]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[23]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[23]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[23]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[23]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[24]~FF  (.D(n874), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[24]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[24]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[24]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[24]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[24]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[24]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[25]~FF  (.D(n872), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[25]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[25]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[25]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[25]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[25]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[25]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[26]~FF  (.D(n870), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[26]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[26]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[26]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[26]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[26]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[26]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[27]~FF  (.D(n868), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[27]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[27]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[27]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[27]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[27]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[27]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[28]~FF  (.D(n866), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[28]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[28]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[28]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[28]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[28]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[28]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[29]~FF  (.D(n864), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[29]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[29]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[29]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[29]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[29]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[29]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[30]~FF  (.D(n862), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[30]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[30]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[30]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[30]~FF .D_POLARITY = 1'b0;
    defparam \useone/H7[30]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[30]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useone/H7[31]~FF  (.D(n861), .CE(\useone/select_1072/Select_2/n3 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useone/H7[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \useone/H7[31]~FF .CLK_POLARITY = 1'b1;
    defparam \useone/H7[31]~FF .CE_POLARITY = 1'b1;
    defparam \useone/H7[31]~FF .SR_POLARITY = 1'b1;
    defparam \useone/H7[31]~FF .D_POLARITY = 1'b1;
    defparam \useone/H7[31]~FF .SR_SYNC = 1'b1;
    defparam \useone/H7[31]~FF .SR_VALUE = 1'b0;
    defparam \useone/H7[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[1]~FF  (.D(\useone/select_1071/Select_1/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[1]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[1]~FF .CE_POLARITY = 1'b1;
    defparam \signature[1]~FF .SR_POLARITY = 1'b1;
    defparam \signature[1]~FF .D_POLARITY = 1'b1;
    defparam \signature[1]~FF .SR_SYNC = 1'b1;
    defparam \signature[1]~FF .SR_VALUE = 1'b0;
    defparam \signature[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[2]~FF  (.D(\useone/n39297 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\signature[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[2]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[2]~FF .CE_POLARITY = 1'b1;
    defparam \signature[2]~FF .SR_POLARITY = 1'b1;
    defparam \signature[2]~FF .D_POLARITY = 1'b1;
    defparam \signature[2]~FF .SR_SYNC = 1'b1;
    defparam \signature[2]~FF .SR_VALUE = 1'b0;
    defparam \signature[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[3]~FF  (.D(\useone/select_1071/Select_3/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[3]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[3]~FF .CE_POLARITY = 1'b1;
    defparam \signature[3]~FF .SR_POLARITY = 1'b1;
    defparam \signature[3]~FF .D_POLARITY = 1'b1;
    defparam \signature[3]~FF .SR_SYNC = 1'b1;
    defparam \signature[3]~FF .SR_VALUE = 1'b0;
    defparam \signature[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[4]~FF  (.D(\useone/select_1071/Select_4/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[4]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[4]~FF .CE_POLARITY = 1'b1;
    defparam \signature[4]~FF .SR_POLARITY = 1'b1;
    defparam \signature[4]~FF .D_POLARITY = 1'b1;
    defparam \signature[4]~FF .SR_SYNC = 1'b1;
    defparam \signature[4]~FF .SR_VALUE = 1'b0;
    defparam \signature[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[5]~FF  (.D(\useone/select_1071/Select_5/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[5]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[5]~FF .CE_POLARITY = 1'b1;
    defparam \signature[5]~FF .SR_POLARITY = 1'b1;
    defparam \signature[5]~FF .D_POLARITY = 1'b1;
    defparam \signature[5]~FF .SR_SYNC = 1'b1;
    defparam \signature[5]~FF .SR_VALUE = 1'b0;
    defparam \signature[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[6]~FF  (.D(\useone/n39293 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\signature[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[6]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[6]~FF .CE_POLARITY = 1'b1;
    defparam \signature[6]~FF .SR_POLARITY = 1'b1;
    defparam \signature[6]~FF .D_POLARITY = 1'b1;
    defparam \signature[6]~FF .SR_SYNC = 1'b1;
    defparam \signature[6]~FF .SR_VALUE = 1'b0;
    defparam \signature[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[7]~FF  (.D(\useone/select_1071/Select_7/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[7]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[7]~FF .CE_POLARITY = 1'b1;
    defparam \signature[7]~FF .SR_POLARITY = 1'b1;
    defparam \signature[7]~FF .D_POLARITY = 1'b1;
    defparam \signature[7]~FF .SR_SYNC = 1'b1;
    defparam \signature[7]~FF .SR_VALUE = 1'b0;
    defparam \signature[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[8]~FF  (.D(\useone/select_1071/Select_8/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[8]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[8]~FF .CE_POLARITY = 1'b1;
    defparam \signature[8]~FF .SR_POLARITY = 1'b1;
    defparam \signature[8]~FF .D_POLARITY = 1'b1;
    defparam \signature[8]~FF .SR_SYNC = 1'b1;
    defparam \signature[8]~FF .SR_VALUE = 1'b0;
    defparam \signature[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[9]~FF  (.D(\useone/select_1071/Select_9/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[9]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[9]~FF .CE_POLARITY = 1'b1;
    defparam \signature[9]~FF .SR_POLARITY = 1'b1;
    defparam \signature[9]~FF .D_POLARITY = 1'b1;
    defparam \signature[9]~FF .SR_SYNC = 1'b1;
    defparam \signature[9]~FF .SR_VALUE = 1'b0;
    defparam \signature[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[10]~FF  (.D(\useone/select_1071/Select_10/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[10]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[10]~FF .CE_POLARITY = 1'b1;
    defparam \signature[10]~FF .SR_POLARITY = 1'b1;
    defparam \signature[10]~FF .D_POLARITY = 1'b1;
    defparam \signature[10]~FF .SR_SYNC = 1'b1;
    defparam \signature[10]~FF .SR_VALUE = 1'b0;
    defparam \signature[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[11]~FF  (.D(\useone/select_1071/Select_11/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[11]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[11]~FF .CE_POLARITY = 1'b1;
    defparam \signature[11]~FF .SR_POLARITY = 1'b1;
    defparam \signature[11]~FF .D_POLARITY = 1'b1;
    defparam \signature[11]~FF .SR_SYNC = 1'b1;
    defparam \signature[11]~FF .SR_VALUE = 1'b0;
    defparam \signature[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[12]~FF  (.D(\useone/select_1071/Select_12/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[12]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[12]~FF .CE_POLARITY = 1'b1;
    defparam \signature[12]~FF .SR_POLARITY = 1'b1;
    defparam \signature[12]~FF .D_POLARITY = 1'b1;
    defparam \signature[12]~FF .SR_SYNC = 1'b1;
    defparam \signature[12]~FF .SR_VALUE = 1'b0;
    defparam \signature[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[13]~FF  (.D(\useone/select_1071/Select_13/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[13]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[13]~FF .CE_POLARITY = 1'b1;
    defparam \signature[13]~FF .SR_POLARITY = 1'b1;
    defparam \signature[13]~FF .D_POLARITY = 1'b1;
    defparam \signature[13]~FF .SR_SYNC = 1'b1;
    defparam \signature[13]~FF .SR_VALUE = 1'b0;
    defparam \signature[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[14]~FF  (.D(\useone/select_1071/Select_14/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[14]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[14]~FF .CE_POLARITY = 1'b1;
    defparam \signature[14]~FF .SR_POLARITY = 1'b1;
    defparam \signature[14]~FF .D_POLARITY = 1'b1;
    defparam \signature[14]~FF .SR_SYNC = 1'b1;
    defparam \signature[14]~FF .SR_VALUE = 1'b0;
    defparam \signature[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[15]~FF  (.D(\useone/n39284 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\signature[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[15]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[15]~FF .CE_POLARITY = 1'b1;
    defparam \signature[15]~FF .SR_POLARITY = 1'b1;
    defparam \signature[15]~FF .D_POLARITY = 1'b1;
    defparam \signature[15]~FF .SR_SYNC = 1'b1;
    defparam \signature[15]~FF .SR_VALUE = 1'b0;
    defparam \signature[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[16]~FF  (.D(\useone/select_1071/Select_16/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[16]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[16]~FF .CE_POLARITY = 1'b1;
    defparam \signature[16]~FF .SR_POLARITY = 1'b1;
    defparam \signature[16]~FF .D_POLARITY = 1'b1;
    defparam \signature[16]~FF .SR_SYNC = 1'b1;
    defparam \signature[16]~FF .SR_VALUE = 1'b0;
    defparam \signature[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[17]~FF  (.D(\useone/select_1071/Select_17/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[17]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[17]~FF .CE_POLARITY = 1'b1;
    defparam \signature[17]~FF .SR_POLARITY = 1'b1;
    defparam \signature[17]~FF .D_POLARITY = 1'b1;
    defparam \signature[17]~FF .SR_SYNC = 1'b1;
    defparam \signature[17]~FF .SR_VALUE = 1'b0;
    defparam \signature[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[18]~FF  (.D(\useone/select_1071/Select_18/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[18]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[18]~FF .CE_POLARITY = 1'b1;
    defparam \signature[18]~FF .SR_POLARITY = 1'b1;
    defparam \signature[18]~FF .D_POLARITY = 1'b1;
    defparam \signature[18]~FF .SR_SYNC = 1'b1;
    defparam \signature[18]~FF .SR_VALUE = 1'b0;
    defparam \signature[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[19]~FF  (.D(\useone/select_1071/Select_19/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[19]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[19]~FF .CE_POLARITY = 1'b1;
    defparam \signature[19]~FF .SR_POLARITY = 1'b1;
    defparam \signature[19]~FF .D_POLARITY = 1'b1;
    defparam \signature[19]~FF .SR_SYNC = 1'b1;
    defparam \signature[19]~FF .SR_VALUE = 1'b0;
    defparam \signature[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[20]~FF  (.D(\useone/select_1071/Select_20/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[20]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[20]~FF .CE_POLARITY = 1'b1;
    defparam \signature[20]~FF .SR_POLARITY = 1'b1;
    defparam \signature[20]~FF .D_POLARITY = 1'b1;
    defparam \signature[20]~FF .SR_SYNC = 1'b1;
    defparam \signature[20]~FF .SR_VALUE = 1'b0;
    defparam \signature[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[21]~FF  (.D(\useone/select_1071/Select_21/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[21]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[21]~FF .CE_POLARITY = 1'b1;
    defparam \signature[21]~FF .SR_POLARITY = 1'b1;
    defparam \signature[21]~FF .D_POLARITY = 1'b1;
    defparam \signature[21]~FF .SR_SYNC = 1'b1;
    defparam \signature[21]~FF .SR_VALUE = 1'b0;
    defparam \signature[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[22]~FF  (.D(\useone/select_1071/Select_22/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[22]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[22]~FF .CE_POLARITY = 1'b1;
    defparam \signature[22]~FF .SR_POLARITY = 1'b1;
    defparam \signature[22]~FF .D_POLARITY = 1'b1;
    defparam \signature[22]~FF .SR_SYNC = 1'b1;
    defparam \signature[22]~FF .SR_VALUE = 1'b0;
    defparam \signature[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[23]~FF  (.D(\useone/select_1071/Select_23/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[23]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[23]~FF .CE_POLARITY = 1'b1;
    defparam \signature[23]~FF .SR_POLARITY = 1'b1;
    defparam \signature[23]~FF .D_POLARITY = 1'b1;
    defparam \signature[23]~FF .SR_SYNC = 1'b1;
    defparam \signature[23]~FF .SR_VALUE = 1'b0;
    defparam \signature[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[24]~FF  (.D(\useone/select_1071/Select_24/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[24]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[24]~FF .CE_POLARITY = 1'b1;
    defparam \signature[24]~FF .SR_POLARITY = 1'b1;
    defparam \signature[24]~FF .D_POLARITY = 1'b1;
    defparam \signature[24]~FF .SR_SYNC = 1'b1;
    defparam \signature[24]~FF .SR_VALUE = 1'b0;
    defparam \signature[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[25]~FF  (.D(\useone/select_1071/Select_25/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[25]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[25]~FF .CE_POLARITY = 1'b1;
    defparam \signature[25]~FF .SR_POLARITY = 1'b1;
    defparam \signature[25]~FF .D_POLARITY = 1'b1;
    defparam \signature[25]~FF .SR_SYNC = 1'b1;
    defparam \signature[25]~FF .SR_VALUE = 1'b0;
    defparam \signature[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[26]~FF  (.D(\useone/select_1071/Select_26/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[26]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[26]~FF .CE_POLARITY = 1'b1;
    defparam \signature[26]~FF .SR_POLARITY = 1'b1;
    defparam \signature[26]~FF .D_POLARITY = 1'b1;
    defparam \signature[26]~FF .SR_SYNC = 1'b1;
    defparam \signature[26]~FF .SR_VALUE = 1'b0;
    defparam \signature[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[27]~FF  (.D(\useone/select_1071/Select_27/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[27]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[27]~FF .CE_POLARITY = 1'b1;
    defparam \signature[27]~FF .SR_POLARITY = 1'b1;
    defparam \signature[27]~FF .D_POLARITY = 1'b1;
    defparam \signature[27]~FF .SR_SYNC = 1'b1;
    defparam \signature[27]~FF .SR_VALUE = 1'b0;
    defparam \signature[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[28]~FF  (.D(\useone/select_1071/Select_28/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[28]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[28]~FF .CE_POLARITY = 1'b1;
    defparam \signature[28]~FF .SR_POLARITY = 1'b1;
    defparam \signature[28]~FF .D_POLARITY = 1'b1;
    defparam \signature[28]~FF .SR_SYNC = 1'b1;
    defparam \signature[28]~FF .SR_VALUE = 1'b0;
    defparam \signature[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[29]~FF  (.D(\useone/select_1071/Select_29/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[29]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[29]~FF .CE_POLARITY = 1'b1;
    defparam \signature[29]~FF .SR_POLARITY = 1'b1;
    defparam \signature[29]~FF .D_POLARITY = 1'b1;
    defparam \signature[29]~FF .SR_SYNC = 1'b1;
    defparam \signature[29]~FF .SR_VALUE = 1'b0;
    defparam \signature[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[30]~FF  (.D(\useone/select_1071/Select_30/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[30]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[30]~FF .CE_POLARITY = 1'b1;
    defparam \signature[30]~FF .SR_POLARITY = 1'b1;
    defparam \signature[30]~FF .D_POLARITY = 1'b1;
    defparam \signature[30]~FF .SR_SYNC = 1'b1;
    defparam \signature[30]~FF .SR_VALUE = 1'b0;
    defparam \signature[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[31]~FF  (.D(\useone/select_1071/Select_31/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[31]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[31]~FF .CE_POLARITY = 1'b1;
    defparam \signature[31]~FF .SR_POLARITY = 1'b1;
    defparam \signature[31]~FF .D_POLARITY = 1'b1;
    defparam \signature[31]~FF .SR_SYNC = 1'b1;
    defparam \signature[31]~FF .SR_VALUE = 1'b0;
    defparam \signature[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[32]~FF  (.D(\useone/select_1071/Select_32/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[32]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[32]~FF .CE_POLARITY = 1'b1;
    defparam \signature[32]~FF .SR_POLARITY = 1'b1;
    defparam \signature[32]~FF .D_POLARITY = 1'b1;
    defparam \signature[32]~FF .SR_SYNC = 1'b1;
    defparam \signature[32]~FF .SR_VALUE = 1'b0;
    defparam \signature[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[33]~FF  (.D(\useone/select_1071/Select_33/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[33]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[33]~FF .CE_POLARITY = 1'b1;
    defparam \signature[33]~FF .SR_POLARITY = 1'b1;
    defparam \signature[33]~FF .D_POLARITY = 1'b1;
    defparam \signature[33]~FF .SR_SYNC = 1'b1;
    defparam \signature[33]~FF .SR_VALUE = 1'b0;
    defparam \signature[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[34]~FF  (.D(\useone/select_1071/Select_34/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[34]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[34]~FF .CE_POLARITY = 1'b1;
    defparam \signature[34]~FF .SR_POLARITY = 1'b1;
    defparam \signature[34]~FF .D_POLARITY = 1'b1;
    defparam \signature[34]~FF .SR_SYNC = 1'b1;
    defparam \signature[34]~FF .SR_VALUE = 1'b0;
    defparam \signature[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[35]~FF  (.D(\useone/select_1071/Select_35/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[35]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[35]~FF .CE_POLARITY = 1'b1;
    defparam \signature[35]~FF .SR_POLARITY = 1'b1;
    defparam \signature[35]~FF .D_POLARITY = 1'b1;
    defparam \signature[35]~FF .SR_SYNC = 1'b1;
    defparam \signature[35]~FF .SR_VALUE = 1'b0;
    defparam \signature[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[36]~FF  (.D(\useone/select_1071/Select_36/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[36]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[36]~FF .CE_POLARITY = 1'b1;
    defparam \signature[36]~FF .SR_POLARITY = 1'b1;
    defparam \signature[36]~FF .D_POLARITY = 1'b1;
    defparam \signature[36]~FF .SR_SYNC = 1'b1;
    defparam \signature[36]~FF .SR_VALUE = 1'b0;
    defparam \signature[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[37]~FF  (.D(\useone/select_1071/Select_37/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[37]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[37]~FF .CE_POLARITY = 1'b1;
    defparam \signature[37]~FF .SR_POLARITY = 1'b1;
    defparam \signature[37]~FF .D_POLARITY = 1'b1;
    defparam \signature[37]~FF .SR_SYNC = 1'b1;
    defparam \signature[37]~FF .SR_VALUE = 1'b0;
    defparam \signature[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[38]~FF  (.D(\useone/select_1071/Select_38/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[38]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[38]~FF .CE_POLARITY = 1'b1;
    defparam \signature[38]~FF .SR_POLARITY = 1'b1;
    defparam \signature[38]~FF .D_POLARITY = 1'b1;
    defparam \signature[38]~FF .SR_SYNC = 1'b1;
    defparam \signature[38]~FF .SR_VALUE = 1'b0;
    defparam \signature[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[39]~FF  (.D(\useone/select_1071/Select_39/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[39]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[39]~FF .CE_POLARITY = 1'b1;
    defparam \signature[39]~FF .SR_POLARITY = 1'b1;
    defparam \signature[39]~FF .D_POLARITY = 1'b1;
    defparam \signature[39]~FF .SR_SYNC = 1'b1;
    defparam \signature[39]~FF .SR_VALUE = 1'b0;
    defparam \signature[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[40]~FF  (.D(\useone/select_1071/Select_40/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[40]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[40]~FF .CE_POLARITY = 1'b1;
    defparam \signature[40]~FF .SR_POLARITY = 1'b1;
    defparam \signature[40]~FF .D_POLARITY = 1'b1;
    defparam \signature[40]~FF .SR_SYNC = 1'b1;
    defparam \signature[40]~FF .SR_VALUE = 1'b0;
    defparam \signature[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[41]~FF  (.D(\useone/select_1071/Select_41/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[41]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[41]~FF .CE_POLARITY = 1'b1;
    defparam \signature[41]~FF .SR_POLARITY = 1'b1;
    defparam \signature[41]~FF .D_POLARITY = 1'b1;
    defparam \signature[41]~FF .SR_SYNC = 1'b1;
    defparam \signature[41]~FF .SR_VALUE = 1'b0;
    defparam \signature[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[42]~FF  (.D(\useone/select_1071/Select_42/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[42]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[42]~FF .CE_POLARITY = 1'b1;
    defparam \signature[42]~FF .SR_POLARITY = 1'b1;
    defparam \signature[42]~FF .D_POLARITY = 1'b1;
    defparam \signature[42]~FF .SR_SYNC = 1'b1;
    defparam \signature[42]~FF .SR_VALUE = 1'b0;
    defparam \signature[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[43]~FF  (.D(\useone/select_1071/Select_43/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[43]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[43]~FF .CE_POLARITY = 1'b1;
    defparam \signature[43]~FF .SR_POLARITY = 1'b1;
    defparam \signature[43]~FF .D_POLARITY = 1'b1;
    defparam \signature[43]~FF .SR_SYNC = 1'b1;
    defparam \signature[43]~FF .SR_VALUE = 1'b0;
    defparam \signature[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[44]~FF  (.D(\useone/select_1071/Select_44/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[44]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[44]~FF .CE_POLARITY = 1'b1;
    defparam \signature[44]~FF .SR_POLARITY = 1'b1;
    defparam \signature[44]~FF .D_POLARITY = 1'b1;
    defparam \signature[44]~FF .SR_SYNC = 1'b1;
    defparam \signature[44]~FF .SR_VALUE = 1'b0;
    defparam \signature[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[45]~FF  (.D(\useone/select_1071/Select_45/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[45]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[45]~FF .CE_POLARITY = 1'b1;
    defparam \signature[45]~FF .SR_POLARITY = 1'b1;
    defparam \signature[45]~FF .D_POLARITY = 1'b1;
    defparam \signature[45]~FF .SR_SYNC = 1'b1;
    defparam \signature[45]~FF .SR_VALUE = 1'b0;
    defparam \signature[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[46]~FF  (.D(\useone/select_1071/Select_46/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[46]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[46]~FF .CE_POLARITY = 1'b1;
    defparam \signature[46]~FF .SR_POLARITY = 1'b1;
    defparam \signature[46]~FF .D_POLARITY = 1'b1;
    defparam \signature[46]~FF .SR_SYNC = 1'b1;
    defparam \signature[46]~FF .SR_VALUE = 1'b0;
    defparam \signature[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[47]~FF  (.D(\useone/select_1071/Select_47/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[47]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[47]~FF .CE_POLARITY = 1'b1;
    defparam \signature[47]~FF .SR_POLARITY = 1'b1;
    defparam \signature[47]~FF .D_POLARITY = 1'b1;
    defparam \signature[47]~FF .SR_SYNC = 1'b1;
    defparam \signature[47]~FF .SR_VALUE = 1'b0;
    defparam \signature[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[48]~FF  (.D(\useone/select_1071/Select_48/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[48]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[48]~FF .CE_POLARITY = 1'b1;
    defparam \signature[48]~FF .SR_POLARITY = 1'b1;
    defparam \signature[48]~FF .D_POLARITY = 1'b1;
    defparam \signature[48]~FF .SR_SYNC = 1'b1;
    defparam \signature[48]~FF .SR_VALUE = 1'b0;
    defparam \signature[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[49]~FF  (.D(\useone/select_1071/Select_49/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[49]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[49]~FF .CE_POLARITY = 1'b1;
    defparam \signature[49]~FF .SR_POLARITY = 1'b1;
    defparam \signature[49]~FF .D_POLARITY = 1'b1;
    defparam \signature[49]~FF .SR_SYNC = 1'b1;
    defparam \signature[49]~FF .SR_VALUE = 1'b0;
    defparam \signature[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[50]~FF  (.D(\useone/select_1071/Select_50/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[50]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[50]~FF .CE_POLARITY = 1'b1;
    defparam \signature[50]~FF .SR_POLARITY = 1'b1;
    defparam \signature[50]~FF .D_POLARITY = 1'b1;
    defparam \signature[50]~FF .SR_SYNC = 1'b1;
    defparam \signature[50]~FF .SR_VALUE = 1'b0;
    defparam \signature[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[51]~FF  (.D(\useone/select_1071/Select_51/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[51]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[51]~FF .CE_POLARITY = 1'b1;
    defparam \signature[51]~FF .SR_POLARITY = 1'b1;
    defparam \signature[51]~FF .D_POLARITY = 1'b1;
    defparam \signature[51]~FF .SR_SYNC = 1'b1;
    defparam \signature[51]~FF .SR_VALUE = 1'b0;
    defparam \signature[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[52]~FF  (.D(\useone/select_1071/Select_52/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[52]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[52]~FF .CE_POLARITY = 1'b1;
    defparam \signature[52]~FF .SR_POLARITY = 1'b1;
    defparam \signature[52]~FF .D_POLARITY = 1'b1;
    defparam \signature[52]~FF .SR_SYNC = 1'b1;
    defparam \signature[52]~FF .SR_VALUE = 1'b0;
    defparam \signature[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[53]~FF  (.D(\useone/select_1071/Select_53/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[53]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[53]~FF .CE_POLARITY = 1'b1;
    defparam \signature[53]~FF .SR_POLARITY = 1'b1;
    defparam \signature[53]~FF .D_POLARITY = 1'b1;
    defparam \signature[53]~FF .SR_SYNC = 1'b1;
    defparam \signature[53]~FF .SR_VALUE = 1'b0;
    defparam \signature[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[54]~FF  (.D(\useone/select_1071/Select_54/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[54]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[54]~FF .CE_POLARITY = 1'b1;
    defparam \signature[54]~FF .SR_POLARITY = 1'b1;
    defparam \signature[54]~FF .D_POLARITY = 1'b1;
    defparam \signature[54]~FF .SR_SYNC = 1'b1;
    defparam \signature[54]~FF .SR_VALUE = 1'b0;
    defparam \signature[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[55]~FF  (.D(\useone/select_1071/Select_55/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[55]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[55]~FF .CE_POLARITY = 1'b1;
    defparam \signature[55]~FF .SR_POLARITY = 1'b1;
    defparam \signature[55]~FF .D_POLARITY = 1'b1;
    defparam \signature[55]~FF .SR_SYNC = 1'b1;
    defparam \signature[55]~FF .SR_VALUE = 1'b0;
    defparam \signature[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[56]~FF  (.D(\useone/select_1071/Select_56/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[56]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[56]~FF .CE_POLARITY = 1'b1;
    defparam \signature[56]~FF .SR_POLARITY = 1'b1;
    defparam \signature[56]~FF .D_POLARITY = 1'b1;
    defparam \signature[56]~FF .SR_SYNC = 1'b1;
    defparam \signature[56]~FF .SR_VALUE = 1'b0;
    defparam \signature[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[57]~FF  (.D(\useone/select_1071/Select_57/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[57]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[57]~FF .CE_POLARITY = 1'b1;
    defparam \signature[57]~FF .SR_POLARITY = 1'b1;
    defparam \signature[57]~FF .D_POLARITY = 1'b1;
    defparam \signature[57]~FF .SR_SYNC = 1'b1;
    defparam \signature[57]~FF .SR_VALUE = 1'b0;
    defparam \signature[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[58]~FF  (.D(\useone/select_1071/Select_58/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[58]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[58]~FF .CE_POLARITY = 1'b1;
    defparam \signature[58]~FF .SR_POLARITY = 1'b1;
    defparam \signature[58]~FF .D_POLARITY = 1'b1;
    defparam \signature[58]~FF .SR_SYNC = 1'b1;
    defparam \signature[58]~FF .SR_VALUE = 1'b0;
    defparam \signature[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[59]~FF  (.D(\useone/select_1071/Select_59/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[59]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[59]~FF .CE_POLARITY = 1'b1;
    defparam \signature[59]~FF .SR_POLARITY = 1'b1;
    defparam \signature[59]~FF .D_POLARITY = 1'b1;
    defparam \signature[59]~FF .SR_SYNC = 1'b1;
    defparam \signature[59]~FF .SR_VALUE = 1'b0;
    defparam \signature[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[60]~FF  (.D(\useone/n39239 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\signature[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[60]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[60]~FF .CE_POLARITY = 1'b1;
    defparam \signature[60]~FF .SR_POLARITY = 1'b1;
    defparam \signature[60]~FF .D_POLARITY = 1'b1;
    defparam \signature[60]~FF .SR_SYNC = 1'b1;
    defparam \signature[60]~FF .SR_VALUE = 1'b0;
    defparam \signature[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[61]~FF  (.D(\useone/select_1071/Select_61/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[61]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[61]~FF .CE_POLARITY = 1'b1;
    defparam \signature[61]~FF .SR_POLARITY = 1'b1;
    defparam \signature[61]~FF .D_POLARITY = 1'b1;
    defparam \signature[61]~FF .SR_SYNC = 1'b1;
    defparam \signature[61]~FF .SR_VALUE = 1'b0;
    defparam \signature[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[62]~FF  (.D(\useone/select_1071/Select_62/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[62]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[62]~FF .CE_POLARITY = 1'b1;
    defparam \signature[62]~FF .SR_POLARITY = 1'b1;
    defparam \signature[62]~FF .D_POLARITY = 1'b1;
    defparam \signature[62]~FF .SR_SYNC = 1'b1;
    defparam \signature[62]~FF .SR_VALUE = 1'b0;
    defparam \signature[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[63]~FF  (.D(\useone/select_1071/Select_63/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[63]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[63]~FF .CE_POLARITY = 1'b1;
    defparam \signature[63]~FF .SR_POLARITY = 1'b1;
    defparam \signature[63]~FF .D_POLARITY = 1'b1;
    defparam \signature[63]~FF .SR_SYNC = 1'b1;
    defparam \signature[63]~FF .SR_VALUE = 1'b0;
    defparam \signature[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[64]~FF  (.D(\useone/select_1071/Select_64/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[64]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[64]~FF .CE_POLARITY = 1'b1;
    defparam \signature[64]~FF .SR_POLARITY = 1'b1;
    defparam \signature[64]~FF .D_POLARITY = 1'b1;
    defparam \signature[64]~FF .SR_SYNC = 1'b1;
    defparam \signature[64]~FF .SR_VALUE = 1'b0;
    defparam \signature[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[65]~FF  (.D(\useone/select_1071/Select_65/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[65]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[65]~FF .CE_POLARITY = 1'b1;
    defparam \signature[65]~FF .SR_POLARITY = 1'b1;
    defparam \signature[65]~FF .D_POLARITY = 1'b1;
    defparam \signature[65]~FF .SR_SYNC = 1'b1;
    defparam \signature[65]~FF .SR_VALUE = 1'b0;
    defparam \signature[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[66]~FF  (.D(\useone/select_1071/Select_66/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[66]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[66]~FF .CE_POLARITY = 1'b1;
    defparam \signature[66]~FF .SR_POLARITY = 1'b1;
    defparam \signature[66]~FF .D_POLARITY = 1'b1;
    defparam \signature[66]~FF .SR_SYNC = 1'b1;
    defparam \signature[66]~FF .SR_VALUE = 1'b0;
    defparam \signature[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[67]~FF  (.D(\useone/select_1071/Select_67/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[67]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[67]~FF .CE_POLARITY = 1'b1;
    defparam \signature[67]~FF .SR_POLARITY = 1'b1;
    defparam \signature[67]~FF .D_POLARITY = 1'b1;
    defparam \signature[67]~FF .SR_SYNC = 1'b1;
    defparam \signature[67]~FF .SR_VALUE = 1'b0;
    defparam \signature[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[68]~FF  (.D(\useone/select_1071/Select_68/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[68]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[68]~FF .CE_POLARITY = 1'b1;
    defparam \signature[68]~FF .SR_POLARITY = 1'b1;
    defparam \signature[68]~FF .D_POLARITY = 1'b1;
    defparam \signature[68]~FF .SR_SYNC = 1'b1;
    defparam \signature[68]~FF .SR_VALUE = 1'b0;
    defparam \signature[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[69]~FF  (.D(\useone/select_1071/Select_69/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[69]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[69]~FF .CE_POLARITY = 1'b1;
    defparam \signature[69]~FF .SR_POLARITY = 1'b1;
    defparam \signature[69]~FF .D_POLARITY = 1'b1;
    defparam \signature[69]~FF .SR_SYNC = 1'b1;
    defparam \signature[69]~FF .SR_VALUE = 1'b0;
    defparam \signature[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[70]~FF  (.D(\useone/select_1071/Select_70/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[70]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[70]~FF .CE_POLARITY = 1'b1;
    defparam \signature[70]~FF .SR_POLARITY = 1'b1;
    defparam \signature[70]~FF .D_POLARITY = 1'b1;
    defparam \signature[70]~FF .SR_SYNC = 1'b1;
    defparam \signature[70]~FF .SR_VALUE = 1'b0;
    defparam \signature[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[71]~FF  (.D(\useone/select_1071/Select_71/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[71]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[71]~FF .CE_POLARITY = 1'b1;
    defparam \signature[71]~FF .SR_POLARITY = 1'b1;
    defparam \signature[71]~FF .D_POLARITY = 1'b1;
    defparam \signature[71]~FF .SR_SYNC = 1'b1;
    defparam \signature[71]~FF .SR_VALUE = 1'b0;
    defparam \signature[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[72]~FF  (.D(\useone/select_1071/Select_72/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[72]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[72]~FF .CE_POLARITY = 1'b1;
    defparam \signature[72]~FF .SR_POLARITY = 1'b1;
    defparam \signature[72]~FF .D_POLARITY = 1'b1;
    defparam \signature[72]~FF .SR_SYNC = 1'b1;
    defparam \signature[72]~FF .SR_VALUE = 1'b0;
    defparam \signature[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[73]~FF  (.D(\useone/select_1071/Select_73/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[73]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[73]~FF .CE_POLARITY = 1'b1;
    defparam \signature[73]~FF .SR_POLARITY = 1'b1;
    defparam \signature[73]~FF .D_POLARITY = 1'b1;
    defparam \signature[73]~FF .SR_SYNC = 1'b1;
    defparam \signature[73]~FF .SR_VALUE = 1'b0;
    defparam \signature[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[74]~FF  (.D(\useone/select_1071/Select_74/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[74]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[74]~FF .CE_POLARITY = 1'b1;
    defparam \signature[74]~FF .SR_POLARITY = 1'b1;
    defparam \signature[74]~FF .D_POLARITY = 1'b1;
    defparam \signature[74]~FF .SR_SYNC = 1'b1;
    defparam \signature[74]~FF .SR_VALUE = 1'b0;
    defparam \signature[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[75]~FF  (.D(\useone/select_1071/Select_75/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[75]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[75]~FF .CE_POLARITY = 1'b1;
    defparam \signature[75]~FF .SR_POLARITY = 1'b1;
    defparam \signature[75]~FF .D_POLARITY = 1'b1;
    defparam \signature[75]~FF .SR_SYNC = 1'b1;
    defparam \signature[75]~FF .SR_VALUE = 1'b0;
    defparam \signature[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[76]~FF  (.D(\useone/select_1071/Select_76/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[76]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[76]~FF .CE_POLARITY = 1'b1;
    defparam \signature[76]~FF .SR_POLARITY = 1'b1;
    defparam \signature[76]~FF .D_POLARITY = 1'b1;
    defparam \signature[76]~FF .SR_SYNC = 1'b1;
    defparam \signature[76]~FF .SR_VALUE = 1'b0;
    defparam \signature[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[77]~FF  (.D(\useone/select_1071/Select_77/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[77]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[77]~FF .CE_POLARITY = 1'b1;
    defparam \signature[77]~FF .SR_POLARITY = 1'b1;
    defparam \signature[77]~FF .D_POLARITY = 1'b1;
    defparam \signature[77]~FF .SR_SYNC = 1'b1;
    defparam \signature[77]~FF .SR_VALUE = 1'b0;
    defparam \signature[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[78]~FF  (.D(\useone/select_1071/Select_78/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[78]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[78]~FF .CE_POLARITY = 1'b1;
    defparam \signature[78]~FF .SR_POLARITY = 1'b1;
    defparam \signature[78]~FF .D_POLARITY = 1'b1;
    defparam \signature[78]~FF .SR_SYNC = 1'b1;
    defparam \signature[78]~FF .SR_VALUE = 1'b0;
    defparam \signature[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[79]~FF  (.D(\useone/select_1071/Select_79/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[79]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[79]~FF .CE_POLARITY = 1'b1;
    defparam \signature[79]~FF .SR_POLARITY = 1'b1;
    defparam \signature[79]~FF .D_POLARITY = 1'b1;
    defparam \signature[79]~FF .SR_SYNC = 1'b1;
    defparam \signature[79]~FF .SR_VALUE = 1'b0;
    defparam \signature[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[80]~FF  (.D(\useone/select_1071/Select_80/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[80]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[80]~FF .CE_POLARITY = 1'b1;
    defparam \signature[80]~FF .SR_POLARITY = 1'b1;
    defparam \signature[80]~FF .D_POLARITY = 1'b1;
    defparam \signature[80]~FF .SR_SYNC = 1'b1;
    defparam \signature[80]~FF .SR_VALUE = 1'b0;
    defparam \signature[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[81]~FF  (.D(\useone/select_1071/Select_81/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[81]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[81]~FF .CE_POLARITY = 1'b1;
    defparam \signature[81]~FF .SR_POLARITY = 1'b1;
    defparam \signature[81]~FF .D_POLARITY = 1'b1;
    defparam \signature[81]~FF .SR_SYNC = 1'b1;
    defparam \signature[81]~FF .SR_VALUE = 1'b0;
    defparam \signature[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[82]~FF  (.D(\useone/select_1071/Select_82/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[82]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[82]~FF .CE_POLARITY = 1'b1;
    defparam \signature[82]~FF .SR_POLARITY = 1'b1;
    defparam \signature[82]~FF .D_POLARITY = 1'b1;
    defparam \signature[82]~FF .SR_SYNC = 1'b1;
    defparam \signature[82]~FF .SR_VALUE = 1'b0;
    defparam \signature[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[83]~FF  (.D(\useone/select_1071/Select_83/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[83]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[83]~FF .CE_POLARITY = 1'b1;
    defparam \signature[83]~FF .SR_POLARITY = 1'b1;
    defparam \signature[83]~FF .D_POLARITY = 1'b1;
    defparam \signature[83]~FF .SR_SYNC = 1'b1;
    defparam \signature[83]~FF .SR_VALUE = 1'b0;
    defparam \signature[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[84]~FF  (.D(\useone/select_1071/Select_84/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[84]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[84]~FF .CE_POLARITY = 1'b1;
    defparam \signature[84]~FF .SR_POLARITY = 1'b1;
    defparam \signature[84]~FF .D_POLARITY = 1'b1;
    defparam \signature[84]~FF .SR_SYNC = 1'b1;
    defparam \signature[84]~FF .SR_VALUE = 1'b0;
    defparam \signature[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[85]~FF  (.D(\useone/select_1071/Select_85/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[85]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[85]~FF .CE_POLARITY = 1'b1;
    defparam \signature[85]~FF .SR_POLARITY = 1'b1;
    defparam \signature[85]~FF .D_POLARITY = 1'b1;
    defparam \signature[85]~FF .SR_SYNC = 1'b1;
    defparam \signature[85]~FF .SR_VALUE = 1'b0;
    defparam \signature[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[86]~FF  (.D(\useone/select_1071/Select_86/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[86]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[86]~FF .CE_POLARITY = 1'b1;
    defparam \signature[86]~FF .SR_POLARITY = 1'b1;
    defparam \signature[86]~FF .D_POLARITY = 1'b1;
    defparam \signature[86]~FF .SR_SYNC = 1'b1;
    defparam \signature[86]~FF .SR_VALUE = 1'b0;
    defparam \signature[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[87]~FF  (.D(\useone/select_1071/Select_87/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[87]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[87]~FF .CE_POLARITY = 1'b1;
    defparam \signature[87]~FF .SR_POLARITY = 1'b1;
    defparam \signature[87]~FF .D_POLARITY = 1'b1;
    defparam \signature[87]~FF .SR_SYNC = 1'b1;
    defparam \signature[87]~FF .SR_VALUE = 1'b0;
    defparam \signature[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[88]~FF  (.D(\useone/select_1071/Select_88/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[88]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[88]~FF .CE_POLARITY = 1'b1;
    defparam \signature[88]~FF .SR_POLARITY = 1'b1;
    defparam \signature[88]~FF .D_POLARITY = 1'b1;
    defparam \signature[88]~FF .SR_SYNC = 1'b1;
    defparam \signature[88]~FF .SR_VALUE = 1'b0;
    defparam \signature[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[89]~FF  (.D(\useone/select_1071/Select_89/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[89]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[89]~FF .CE_POLARITY = 1'b1;
    defparam \signature[89]~FF .SR_POLARITY = 1'b1;
    defparam \signature[89]~FF .D_POLARITY = 1'b1;
    defparam \signature[89]~FF .SR_SYNC = 1'b1;
    defparam \signature[89]~FF .SR_VALUE = 1'b0;
    defparam \signature[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[90]~FF  (.D(\useone/select_1071/Select_90/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[90]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[90]~FF .CE_POLARITY = 1'b1;
    defparam \signature[90]~FF .SR_POLARITY = 1'b1;
    defparam \signature[90]~FF .D_POLARITY = 1'b1;
    defparam \signature[90]~FF .SR_SYNC = 1'b1;
    defparam \signature[90]~FF .SR_VALUE = 1'b0;
    defparam \signature[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[91]~FF  (.D(\useone/select_1071/Select_91/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[91]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[91]~FF .CE_POLARITY = 1'b1;
    defparam \signature[91]~FF .SR_POLARITY = 1'b1;
    defparam \signature[91]~FF .D_POLARITY = 1'b1;
    defparam \signature[91]~FF .SR_SYNC = 1'b1;
    defparam \signature[91]~FF .SR_VALUE = 1'b0;
    defparam \signature[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[92]~FF  (.D(\useone/select_1071/Select_92/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[92]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[92]~FF .CE_POLARITY = 1'b1;
    defparam \signature[92]~FF .SR_POLARITY = 1'b1;
    defparam \signature[92]~FF .D_POLARITY = 1'b1;
    defparam \signature[92]~FF .SR_SYNC = 1'b1;
    defparam \signature[92]~FF .SR_VALUE = 1'b0;
    defparam \signature[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[93]~FF  (.D(\useone/select_1071/Select_93/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[93]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[93]~FF .CE_POLARITY = 1'b1;
    defparam \signature[93]~FF .SR_POLARITY = 1'b1;
    defparam \signature[93]~FF .D_POLARITY = 1'b1;
    defparam \signature[93]~FF .SR_SYNC = 1'b1;
    defparam \signature[93]~FF .SR_VALUE = 1'b0;
    defparam \signature[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[94]~FF  (.D(\useone/select_1071/Select_94/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[94]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[94]~FF .CE_POLARITY = 1'b1;
    defparam \signature[94]~FF .SR_POLARITY = 1'b1;
    defparam \signature[94]~FF .D_POLARITY = 1'b1;
    defparam \signature[94]~FF .SR_SYNC = 1'b1;
    defparam \signature[94]~FF .SR_VALUE = 1'b0;
    defparam \signature[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[95]~FF  (.D(\useone/select_1071/Select_95/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[95]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[95]~FF .CE_POLARITY = 1'b1;
    defparam \signature[95]~FF .SR_POLARITY = 1'b1;
    defparam \signature[95]~FF .D_POLARITY = 1'b1;
    defparam \signature[95]~FF .SR_SYNC = 1'b1;
    defparam \signature[95]~FF .SR_VALUE = 1'b0;
    defparam \signature[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[96]~FF  (.D(\useone/select_1071/Select_96/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[96]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[96]~FF .CE_POLARITY = 1'b1;
    defparam \signature[96]~FF .SR_POLARITY = 1'b1;
    defparam \signature[96]~FF .D_POLARITY = 1'b1;
    defparam \signature[96]~FF .SR_SYNC = 1'b1;
    defparam \signature[96]~FF .SR_VALUE = 1'b0;
    defparam \signature[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[97]~FF  (.D(\useone/select_1071/Select_97/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[97]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[97]~FF .CE_POLARITY = 1'b1;
    defparam \signature[97]~FF .SR_POLARITY = 1'b1;
    defparam \signature[97]~FF .D_POLARITY = 1'b1;
    defparam \signature[97]~FF .SR_SYNC = 1'b1;
    defparam \signature[97]~FF .SR_VALUE = 1'b0;
    defparam \signature[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[98]~FF  (.D(\useone/select_1071/Select_98/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[98]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[98]~FF .CE_POLARITY = 1'b1;
    defparam \signature[98]~FF .SR_POLARITY = 1'b1;
    defparam \signature[98]~FF .D_POLARITY = 1'b1;
    defparam \signature[98]~FF .SR_SYNC = 1'b1;
    defparam \signature[98]~FF .SR_VALUE = 1'b0;
    defparam \signature[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[99]~FF  (.D(\useone/select_1071/Select_99/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[99]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[99]~FF .CE_POLARITY = 1'b1;
    defparam \signature[99]~FF .SR_POLARITY = 1'b1;
    defparam \signature[99]~FF .D_POLARITY = 1'b1;
    defparam \signature[99]~FF .SR_SYNC = 1'b1;
    defparam \signature[99]~FF .SR_VALUE = 1'b0;
    defparam \signature[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[100]~FF  (.D(\useone/select_1071/Select_100/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[100]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[100]~FF .CE_POLARITY = 1'b1;
    defparam \signature[100]~FF .SR_POLARITY = 1'b1;
    defparam \signature[100]~FF .D_POLARITY = 1'b1;
    defparam \signature[100]~FF .SR_SYNC = 1'b1;
    defparam \signature[100]~FF .SR_VALUE = 1'b0;
    defparam \signature[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[101]~FF  (.D(\useone/select_1071/Select_101/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[101]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[101]~FF .CE_POLARITY = 1'b1;
    defparam \signature[101]~FF .SR_POLARITY = 1'b1;
    defparam \signature[101]~FF .D_POLARITY = 1'b1;
    defparam \signature[101]~FF .SR_SYNC = 1'b1;
    defparam \signature[101]~FF .SR_VALUE = 1'b0;
    defparam \signature[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[102]~FF  (.D(\useone/select_1071/Select_102/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[102]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[102]~FF .CE_POLARITY = 1'b1;
    defparam \signature[102]~FF .SR_POLARITY = 1'b1;
    defparam \signature[102]~FF .D_POLARITY = 1'b1;
    defparam \signature[102]~FF .SR_SYNC = 1'b1;
    defparam \signature[102]~FF .SR_VALUE = 1'b0;
    defparam \signature[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[103]~FF  (.D(\useone/select_1071/Select_103/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[103]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[103]~FF .CE_POLARITY = 1'b1;
    defparam \signature[103]~FF .SR_POLARITY = 1'b1;
    defparam \signature[103]~FF .D_POLARITY = 1'b1;
    defparam \signature[103]~FF .SR_SYNC = 1'b1;
    defparam \signature[103]~FF .SR_VALUE = 1'b0;
    defparam \signature[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[104]~FF  (.D(\useone/select_1071/Select_104/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[104]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[104]~FF .CE_POLARITY = 1'b1;
    defparam \signature[104]~FF .SR_POLARITY = 1'b1;
    defparam \signature[104]~FF .D_POLARITY = 1'b1;
    defparam \signature[104]~FF .SR_SYNC = 1'b1;
    defparam \signature[104]~FF .SR_VALUE = 1'b0;
    defparam \signature[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[105]~FF  (.D(\useone/select_1071/Select_105/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[105]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[105]~FF .CE_POLARITY = 1'b1;
    defparam \signature[105]~FF .SR_POLARITY = 1'b1;
    defparam \signature[105]~FF .D_POLARITY = 1'b1;
    defparam \signature[105]~FF .SR_SYNC = 1'b1;
    defparam \signature[105]~FF .SR_VALUE = 1'b0;
    defparam \signature[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[106]~FF  (.D(\useone/select_1071/Select_106/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[106]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[106]~FF .CE_POLARITY = 1'b1;
    defparam \signature[106]~FF .SR_POLARITY = 1'b1;
    defparam \signature[106]~FF .D_POLARITY = 1'b1;
    defparam \signature[106]~FF .SR_SYNC = 1'b1;
    defparam \signature[106]~FF .SR_VALUE = 1'b0;
    defparam \signature[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[107]~FF  (.D(\useone/select_1071/Select_107/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[107]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[107]~FF .CE_POLARITY = 1'b1;
    defparam \signature[107]~FF .SR_POLARITY = 1'b1;
    defparam \signature[107]~FF .D_POLARITY = 1'b1;
    defparam \signature[107]~FF .SR_SYNC = 1'b1;
    defparam \signature[107]~FF .SR_VALUE = 1'b0;
    defparam \signature[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[108]~FF  (.D(\useone/select_1071/Select_108/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[108]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[108]~FF .CE_POLARITY = 1'b1;
    defparam \signature[108]~FF .SR_POLARITY = 1'b1;
    defparam \signature[108]~FF .D_POLARITY = 1'b1;
    defparam \signature[108]~FF .SR_SYNC = 1'b1;
    defparam \signature[108]~FF .SR_VALUE = 1'b0;
    defparam \signature[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[109]~FF  (.D(\useone/select_1071/Select_109/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[109]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[109]~FF .CE_POLARITY = 1'b1;
    defparam \signature[109]~FF .SR_POLARITY = 1'b1;
    defparam \signature[109]~FF .D_POLARITY = 1'b1;
    defparam \signature[109]~FF .SR_SYNC = 1'b1;
    defparam \signature[109]~FF .SR_VALUE = 1'b0;
    defparam \signature[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[110]~FF  (.D(\useone/select_1071/Select_110/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[110]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[110]~FF .CE_POLARITY = 1'b1;
    defparam \signature[110]~FF .SR_POLARITY = 1'b1;
    defparam \signature[110]~FF .D_POLARITY = 1'b1;
    defparam \signature[110]~FF .SR_SYNC = 1'b1;
    defparam \signature[110]~FF .SR_VALUE = 1'b0;
    defparam \signature[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[111]~FF  (.D(\useone/select_1071/Select_111/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[111]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[111]~FF .CE_POLARITY = 1'b1;
    defparam \signature[111]~FF .SR_POLARITY = 1'b1;
    defparam \signature[111]~FF .D_POLARITY = 1'b1;
    defparam \signature[111]~FF .SR_SYNC = 1'b1;
    defparam \signature[111]~FF .SR_VALUE = 1'b0;
    defparam \signature[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[112]~FF  (.D(\useone/select_1071/Select_112/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[112]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[112]~FF .CE_POLARITY = 1'b1;
    defparam \signature[112]~FF .SR_POLARITY = 1'b1;
    defparam \signature[112]~FF .D_POLARITY = 1'b1;
    defparam \signature[112]~FF .SR_SYNC = 1'b1;
    defparam \signature[112]~FF .SR_VALUE = 1'b0;
    defparam \signature[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[113]~FF  (.D(\useone/select_1071/Select_113/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[113]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[113]~FF .CE_POLARITY = 1'b1;
    defparam \signature[113]~FF .SR_POLARITY = 1'b1;
    defparam \signature[113]~FF .D_POLARITY = 1'b1;
    defparam \signature[113]~FF .SR_SYNC = 1'b1;
    defparam \signature[113]~FF .SR_VALUE = 1'b0;
    defparam \signature[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[114]~FF  (.D(\useone/select_1071/Select_114/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[114]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[114]~FF .CE_POLARITY = 1'b1;
    defparam \signature[114]~FF .SR_POLARITY = 1'b1;
    defparam \signature[114]~FF .D_POLARITY = 1'b1;
    defparam \signature[114]~FF .SR_SYNC = 1'b1;
    defparam \signature[114]~FF .SR_VALUE = 1'b0;
    defparam \signature[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[115]~FF  (.D(\useone/select_1071/Select_115/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[115]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[115]~FF .CE_POLARITY = 1'b1;
    defparam \signature[115]~FF .SR_POLARITY = 1'b1;
    defparam \signature[115]~FF .D_POLARITY = 1'b1;
    defparam \signature[115]~FF .SR_SYNC = 1'b1;
    defparam \signature[115]~FF .SR_VALUE = 1'b0;
    defparam \signature[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[116]~FF  (.D(\useone/select_1071/Select_116/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[116]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[116]~FF .CE_POLARITY = 1'b1;
    defparam \signature[116]~FF .SR_POLARITY = 1'b1;
    defparam \signature[116]~FF .D_POLARITY = 1'b1;
    defparam \signature[116]~FF .SR_SYNC = 1'b1;
    defparam \signature[116]~FF .SR_VALUE = 1'b0;
    defparam \signature[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[117]~FF  (.D(\useone/select_1071/Select_117/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[117]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[117]~FF .CE_POLARITY = 1'b1;
    defparam \signature[117]~FF .SR_POLARITY = 1'b1;
    defparam \signature[117]~FF .D_POLARITY = 1'b1;
    defparam \signature[117]~FF .SR_SYNC = 1'b1;
    defparam \signature[117]~FF .SR_VALUE = 1'b0;
    defparam \signature[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[118]~FF  (.D(\useone/select_1071/Select_118/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[118]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[118]~FF .CE_POLARITY = 1'b1;
    defparam \signature[118]~FF .SR_POLARITY = 1'b1;
    defparam \signature[118]~FF .D_POLARITY = 1'b1;
    defparam \signature[118]~FF .SR_SYNC = 1'b1;
    defparam \signature[118]~FF .SR_VALUE = 1'b0;
    defparam \signature[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[119]~FF  (.D(\useone/select_1071/Select_119/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[119]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[119]~FF .CE_POLARITY = 1'b1;
    defparam \signature[119]~FF .SR_POLARITY = 1'b1;
    defparam \signature[119]~FF .D_POLARITY = 1'b1;
    defparam \signature[119]~FF .SR_SYNC = 1'b1;
    defparam \signature[119]~FF .SR_VALUE = 1'b0;
    defparam \signature[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[120]~FF  (.D(\useone/select_1071/Select_120/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[120]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[120]~FF .CE_POLARITY = 1'b1;
    defparam \signature[120]~FF .SR_POLARITY = 1'b1;
    defparam \signature[120]~FF .D_POLARITY = 1'b1;
    defparam \signature[120]~FF .SR_SYNC = 1'b1;
    defparam \signature[120]~FF .SR_VALUE = 1'b0;
    defparam \signature[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[121]~FF  (.D(\useone/select_1071/Select_121/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[121]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[121]~FF .CE_POLARITY = 1'b1;
    defparam \signature[121]~FF .SR_POLARITY = 1'b1;
    defparam \signature[121]~FF .D_POLARITY = 1'b1;
    defparam \signature[121]~FF .SR_SYNC = 1'b1;
    defparam \signature[121]~FF .SR_VALUE = 1'b0;
    defparam \signature[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[122]~FF  (.D(\useone/select_1071/Select_122/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[122]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[122]~FF .CE_POLARITY = 1'b1;
    defparam \signature[122]~FF .SR_POLARITY = 1'b1;
    defparam \signature[122]~FF .D_POLARITY = 1'b1;
    defparam \signature[122]~FF .SR_SYNC = 1'b1;
    defparam \signature[122]~FF .SR_VALUE = 1'b0;
    defparam \signature[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[123]~FF  (.D(\useone/select_1071/Select_123/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[123]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[123]~FF .CE_POLARITY = 1'b1;
    defparam \signature[123]~FF .SR_POLARITY = 1'b1;
    defparam \signature[123]~FF .D_POLARITY = 1'b1;
    defparam \signature[123]~FF .SR_SYNC = 1'b1;
    defparam \signature[123]~FF .SR_VALUE = 1'b0;
    defparam \signature[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[124]~FF  (.D(\useone/select_1071/Select_124/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[124]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[124]~FF .CE_POLARITY = 1'b1;
    defparam \signature[124]~FF .SR_POLARITY = 1'b1;
    defparam \signature[124]~FF .D_POLARITY = 1'b1;
    defparam \signature[124]~FF .SR_SYNC = 1'b1;
    defparam \signature[124]~FF .SR_VALUE = 1'b0;
    defparam \signature[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[125]~FF  (.D(\useone/select_1071/Select_125/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[125]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[125]~FF .CE_POLARITY = 1'b1;
    defparam \signature[125]~FF .SR_POLARITY = 1'b1;
    defparam \signature[125]~FF .D_POLARITY = 1'b1;
    defparam \signature[125]~FF .SR_SYNC = 1'b1;
    defparam \signature[125]~FF .SR_VALUE = 1'b0;
    defparam \signature[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[126]~FF  (.D(\useone/select_1071/Select_126/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[126]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[126]~FF .CE_POLARITY = 1'b1;
    defparam \signature[126]~FF .SR_POLARITY = 1'b1;
    defparam \signature[126]~FF .D_POLARITY = 1'b1;
    defparam \signature[126]~FF .SR_SYNC = 1'b1;
    defparam \signature[126]~FF .SR_VALUE = 1'b0;
    defparam \signature[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[127]~FF  (.D(\useone/select_1071/Select_127/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[127]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[127]~FF .CE_POLARITY = 1'b1;
    defparam \signature[127]~FF .SR_POLARITY = 1'b1;
    defparam \signature[127]~FF .D_POLARITY = 1'b1;
    defparam \signature[127]~FF .SR_SYNC = 1'b1;
    defparam \signature[127]~FF .SR_VALUE = 1'b0;
    defparam \signature[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[128]~FF  (.D(\useone/n39171 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\signature[128] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[128]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[128]~FF .CE_POLARITY = 1'b1;
    defparam \signature[128]~FF .SR_POLARITY = 1'b1;
    defparam \signature[128]~FF .D_POLARITY = 1'b1;
    defparam \signature[128]~FF .SR_SYNC = 1'b1;
    defparam \signature[128]~FF .SR_VALUE = 1'b0;
    defparam \signature[128]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[129]~FF  (.D(\useone/select_1071/Select_129/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[129] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[129]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[129]~FF .CE_POLARITY = 1'b1;
    defparam \signature[129]~FF .SR_POLARITY = 1'b1;
    defparam \signature[129]~FF .D_POLARITY = 1'b1;
    defparam \signature[129]~FF .SR_SYNC = 1'b1;
    defparam \signature[129]~FF .SR_VALUE = 1'b0;
    defparam \signature[129]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[130]~FF  (.D(\useone/select_1071/Select_130/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[130] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[130]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[130]~FF .CE_POLARITY = 1'b1;
    defparam \signature[130]~FF .SR_POLARITY = 1'b1;
    defparam \signature[130]~FF .D_POLARITY = 1'b1;
    defparam \signature[130]~FF .SR_SYNC = 1'b1;
    defparam \signature[130]~FF .SR_VALUE = 1'b0;
    defparam \signature[130]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[131]~FF  (.D(\useone/select_1071/Select_131/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[131] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[131]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[131]~FF .CE_POLARITY = 1'b1;
    defparam \signature[131]~FF .SR_POLARITY = 1'b1;
    defparam \signature[131]~FF .D_POLARITY = 1'b1;
    defparam \signature[131]~FF .SR_SYNC = 1'b1;
    defparam \signature[131]~FF .SR_VALUE = 1'b0;
    defparam \signature[131]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[132]~FF  (.D(\useone/n39167 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(1'b0), .Q(\signature[132] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[132]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[132]~FF .CE_POLARITY = 1'b1;
    defparam \signature[132]~FF .SR_POLARITY = 1'b1;
    defparam \signature[132]~FF .D_POLARITY = 1'b1;
    defparam \signature[132]~FF .SR_SYNC = 1'b1;
    defparam \signature[132]~FF .SR_VALUE = 1'b0;
    defparam \signature[132]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[133]~FF  (.D(\useone/select_1071/Select_133/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[133] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[133]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[133]~FF .CE_POLARITY = 1'b1;
    defparam \signature[133]~FF .SR_POLARITY = 1'b1;
    defparam \signature[133]~FF .D_POLARITY = 1'b1;
    defparam \signature[133]~FF .SR_SYNC = 1'b1;
    defparam \signature[133]~FF .SR_VALUE = 1'b0;
    defparam \signature[133]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[134]~FF  (.D(\useone/select_1071/Select_134/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[134] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[134]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[134]~FF .CE_POLARITY = 1'b1;
    defparam \signature[134]~FF .SR_POLARITY = 1'b1;
    defparam \signature[134]~FF .D_POLARITY = 1'b1;
    defparam \signature[134]~FF .SR_SYNC = 1'b1;
    defparam \signature[134]~FF .SR_VALUE = 1'b0;
    defparam \signature[134]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[135]~FF  (.D(\useone/select_1071/Select_135/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[135] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[135]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[135]~FF .CE_POLARITY = 1'b1;
    defparam \signature[135]~FF .SR_POLARITY = 1'b1;
    defparam \signature[135]~FF .D_POLARITY = 1'b1;
    defparam \signature[135]~FF .SR_SYNC = 1'b1;
    defparam \signature[135]~FF .SR_VALUE = 1'b0;
    defparam \signature[135]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[136]~FF  (.D(\useone/select_1071/Select_136/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[136] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[136]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[136]~FF .CE_POLARITY = 1'b1;
    defparam \signature[136]~FF .SR_POLARITY = 1'b1;
    defparam \signature[136]~FF .D_POLARITY = 1'b1;
    defparam \signature[136]~FF .SR_SYNC = 1'b1;
    defparam \signature[136]~FF .SR_VALUE = 1'b0;
    defparam \signature[136]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[137]~FF  (.D(\useone/select_1071/Select_137/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[137] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[137]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[137]~FF .CE_POLARITY = 1'b1;
    defparam \signature[137]~FF .SR_POLARITY = 1'b1;
    defparam \signature[137]~FF .D_POLARITY = 1'b1;
    defparam \signature[137]~FF .SR_SYNC = 1'b1;
    defparam \signature[137]~FF .SR_VALUE = 1'b0;
    defparam \signature[137]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[138]~FF  (.D(\useone/select_1071/Select_138/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[138] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[138]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[138]~FF .CE_POLARITY = 1'b1;
    defparam \signature[138]~FF .SR_POLARITY = 1'b1;
    defparam \signature[138]~FF .D_POLARITY = 1'b1;
    defparam \signature[138]~FF .SR_SYNC = 1'b1;
    defparam \signature[138]~FF .SR_VALUE = 1'b0;
    defparam \signature[138]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[139]~FF  (.D(\useone/select_1071/Select_139/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[139] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[139]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[139]~FF .CE_POLARITY = 1'b1;
    defparam \signature[139]~FF .SR_POLARITY = 1'b1;
    defparam \signature[139]~FF .D_POLARITY = 1'b1;
    defparam \signature[139]~FF .SR_SYNC = 1'b1;
    defparam \signature[139]~FF .SR_VALUE = 1'b0;
    defparam \signature[139]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[140]~FF  (.D(\useone/select_1071/Select_140/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[140] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[140]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[140]~FF .CE_POLARITY = 1'b1;
    defparam \signature[140]~FF .SR_POLARITY = 1'b1;
    defparam \signature[140]~FF .D_POLARITY = 1'b1;
    defparam \signature[140]~FF .SR_SYNC = 1'b1;
    defparam \signature[140]~FF .SR_VALUE = 1'b0;
    defparam \signature[140]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[141]~FF  (.D(\useone/select_1071/Select_141/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[141] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[141]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[141]~FF .CE_POLARITY = 1'b1;
    defparam \signature[141]~FF .SR_POLARITY = 1'b1;
    defparam \signature[141]~FF .D_POLARITY = 1'b1;
    defparam \signature[141]~FF .SR_SYNC = 1'b1;
    defparam \signature[141]~FF .SR_VALUE = 1'b0;
    defparam \signature[141]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[142]~FF  (.D(\useone/select_1071/Select_142/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[142] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[142]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[142]~FF .CE_POLARITY = 1'b1;
    defparam \signature[142]~FF .SR_POLARITY = 1'b1;
    defparam \signature[142]~FF .D_POLARITY = 1'b1;
    defparam \signature[142]~FF .SR_SYNC = 1'b1;
    defparam \signature[142]~FF .SR_VALUE = 1'b0;
    defparam \signature[142]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[143]~FF  (.D(\useone/select_1071/Select_143/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[143] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[143]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[143]~FF .CE_POLARITY = 1'b1;
    defparam \signature[143]~FF .SR_POLARITY = 1'b1;
    defparam \signature[143]~FF .D_POLARITY = 1'b1;
    defparam \signature[143]~FF .SR_SYNC = 1'b1;
    defparam \signature[143]~FF .SR_VALUE = 1'b0;
    defparam \signature[143]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[144]~FF  (.D(\useone/select_1071/Select_144/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[144] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[144]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[144]~FF .CE_POLARITY = 1'b1;
    defparam \signature[144]~FF .SR_POLARITY = 1'b1;
    defparam \signature[144]~FF .D_POLARITY = 1'b1;
    defparam \signature[144]~FF .SR_SYNC = 1'b1;
    defparam \signature[144]~FF .SR_VALUE = 1'b0;
    defparam \signature[144]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[145]~FF  (.D(\useone/select_1071/Select_145/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[145] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[145]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[145]~FF .CE_POLARITY = 1'b1;
    defparam \signature[145]~FF .SR_POLARITY = 1'b1;
    defparam \signature[145]~FF .D_POLARITY = 1'b1;
    defparam \signature[145]~FF .SR_SYNC = 1'b1;
    defparam \signature[145]~FF .SR_VALUE = 1'b0;
    defparam \signature[145]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[146]~FF  (.D(\useone/select_1071/Select_146/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[146] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[146]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[146]~FF .CE_POLARITY = 1'b1;
    defparam \signature[146]~FF .SR_POLARITY = 1'b1;
    defparam \signature[146]~FF .D_POLARITY = 1'b1;
    defparam \signature[146]~FF .SR_SYNC = 1'b1;
    defparam \signature[146]~FF .SR_VALUE = 1'b0;
    defparam \signature[146]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[147]~FF  (.D(\useone/select_1071/Select_147/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[147] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[147]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[147]~FF .CE_POLARITY = 1'b1;
    defparam \signature[147]~FF .SR_POLARITY = 1'b1;
    defparam \signature[147]~FF .D_POLARITY = 1'b1;
    defparam \signature[147]~FF .SR_SYNC = 1'b1;
    defparam \signature[147]~FF .SR_VALUE = 1'b0;
    defparam \signature[147]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[148]~FF  (.D(\useone/select_1071/Select_148/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[148] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[148]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[148]~FF .CE_POLARITY = 1'b1;
    defparam \signature[148]~FF .SR_POLARITY = 1'b1;
    defparam \signature[148]~FF .D_POLARITY = 1'b1;
    defparam \signature[148]~FF .SR_SYNC = 1'b1;
    defparam \signature[148]~FF .SR_VALUE = 1'b0;
    defparam \signature[148]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[149]~FF  (.D(\useone/select_1071/Select_149/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[149] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[149]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[149]~FF .CE_POLARITY = 1'b1;
    defparam \signature[149]~FF .SR_POLARITY = 1'b1;
    defparam \signature[149]~FF .D_POLARITY = 1'b1;
    defparam \signature[149]~FF .SR_SYNC = 1'b1;
    defparam \signature[149]~FF .SR_VALUE = 1'b0;
    defparam \signature[149]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[150]~FF  (.D(\useone/select_1071/Select_150/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[150] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[150]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[150]~FF .CE_POLARITY = 1'b1;
    defparam \signature[150]~FF .SR_POLARITY = 1'b1;
    defparam \signature[150]~FF .D_POLARITY = 1'b1;
    defparam \signature[150]~FF .SR_SYNC = 1'b1;
    defparam \signature[150]~FF .SR_VALUE = 1'b0;
    defparam \signature[150]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[151]~FF  (.D(\useone/select_1071/Select_151/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[151] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[151]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[151]~FF .CE_POLARITY = 1'b1;
    defparam \signature[151]~FF .SR_POLARITY = 1'b1;
    defparam \signature[151]~FF .D_POLARITY = 1'b1;
    defparam \signature[151]~FF .SR_SYNC = 1'b1;
    defparam \signature[151]~FF .SR_VALUE = 1'b0;
    defparam \signature[151]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[152]~FF  (.D(\useone/select_1071/Select_152/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[152] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[152]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[152]~FF .CE_POLARITY = 1'b1;
    defparam \signature[152]~FF .SR_POLARITY = 1'b1;
    defparam \signature[152]~FF .D_POLARITY = 1'b1;
    defparam \signature[152]~FF .SR_SYNC = 1'b1;
    defparam \signature[152]~FF .SR_VALUE = 1'b0;
    defparam \signature[152]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[153]~FF  (.D(\useone/select_1071/Select_153/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[153] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[153]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[153]~FF .CE_POLARITY = 1'b1;
    defparam \signature[153]~FF .SR_POLARITY = 1'b1;
    defparam \signature[153]~FF .D_POLARITY = 1'b1;
    defparam \signature[153]~FF .SR_SYNC = 1'b1;
    defparam \signature[153]~FF .SR_VALUE = 1'b0;
    defparam \signature[153]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[154]~FF  (.D(\useone/select_1071/Select_154/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[154] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[154]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[154]~FF .CE_POLARITY = 1'b1;
    defparam \signature[154]~FF .SR_POLARITY = 1'b1;
    defparam \signature[154]~FF .D_POLARITY = 1'b1;
    defparam \signature[154]~FF .SR_SYNC = 1'b1;
    defparam \signature[154]~FF .SR_VALUE = 1'b0;
    defparam \signature[154]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[155]~FF  (.D(\useone/select_1071/Select_155/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[155] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[155]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[155]~FF .CE_POLARITY = 1'b1;
    defparam \signature[155]~FF .SR_POLARITY = 1'b1;
    defparam \signature[155]~FF .D_POLARITY = 1'b1;
    defparam \signature[155]~FF .SR_SYNC = 1'b1;
    defparam \signature[155]~FF .SR_VALUE = 1'b0;
    defparam \signature[155]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[156]~FF  (.D(\useone/select_1071/Select_156/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[156] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[156]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[156]~FF .CE_POLARITY = 1'b1;
    defparam \signature[156]~FF .SR_POLARITY = 1'b1;
    defparam \signature[156]~FF .D_POLARITY = 1'b1;
    defparam \signature[156]~FF .SR_SYNC = 1'b1;
    defparam \signature[156]~FF .SR_VALUE = 1'b0;
    defparam \signature[156]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[157]~FF  (.D(\useone/select_1071/Select_157/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[157] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[157]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[157]~FF .CE_POLARITY = 1'b1;
    defparam \signature[157]~FF .SR_POLARITY = 1'b1;
    defparam \signature[157]~FF .D_POLARITY = 1'b1;
    defparam \signature[157]~FF .SR_SYNC = 1'b1;
    defparam \signature[157]~FF .SR_VALUE = 1'b0;
    defparam \signature[157]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[158]~FF  (.D(\useone/select_1071/Select_158/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[158] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[158]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[158]~FF .CE_POLARITY = 1'b1;
    defparam \signature[158]~FF .SR_POLARITY = 1'b1;
    defparam \signature[158]~FF .D_POLARITY = 1'b1;
    defparam \signature[158]~FF .SR_SYNC = 1'b1;
    defparam \signature[158]~FF .SR_VALUE = 1'b0;
    defparam \signature[158]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[159]~FF  (.D(\useone/select_1071/Select_159/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[159] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[159]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[159]~FF .CE_POLARITY = 1'b1;
    defparam \signature[159]~FF .SR_POLARITY = 1'b1;
    defparam \signature[159]~FF .D_POLARITY = 1'b1;
    defparam \signature[159]~FF .SR_SYNC = 1'b1;
    defparam \signature[159]~FF .SR_VALUE = 1'b0;
    defparam \signature[159]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[160]~FF  (.D(\useone/select_1071/Select_160/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[160] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[160]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[160]~FF .CE_POLARITY = 1'b1;
    defparam \signature[160]~FF .SR_POLARITY = 1'b1;
    defparam \signature[160]~FF .D_POLARITY = 1'b1;
    defparam \signature[160]~FF .SR_SYNC = 1'b1;
    defparam \signature[160]~FF .SR_VALUE = 1'b0;
    defparam \signature[160]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[161]~FF  (.D(\useone/select_1071/Select_161/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[161] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[161]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[161]~FF .CE_POLARITY = 1'b1;
    defparam \signature[161]~FF .SR_POLARITY = 1'b1;
    defparam \signature[161]~FF .D_POLARITY = 1'b1;
    defparam \signature[161]~FF .SR_SYNC = 1'b1;
    defparam \signature[161]~FF .SR_VALUE = 1'b0;
    defparam \signature[161]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[162]~FF  (.D(\useone/select_1071/Select_162/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[162] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[162]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[162]~FF .CE_POLARITY = 1'b1;
    defparam \signature[162]~FF .SR_POLARITY = 1'b1;
    defparam \signature[162]~FF .D_POLARITY = 1'b1;
    defparam \signature[162]~FF .SR_SYNC = 1'b1;
    defparam \signature[162]~FF .SR_VALUE = 1'b0;
    defparam \signature[162]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[163]~FF  (.D(\useone/select_1071/Select_163/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[163] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[163]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[163]~FF .CE_POLARITY = 1'b1;
    defparam \signature[163]~FF .SR_POLARITY = 1'b1;
    defparam \signature[163]~FF .D_POLARITY = 1'b1;
    defparam \signature[163]~FF .SR_SYNC = 1'b1;
    defparam \signature[163]~FF .SR_VALUE = 1'b0;
    defparam \signature[163]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[164]~FF  (.D(\useone/select_1071/Select_164/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[164] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[164]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[164]~FF .CE_POLARITY = 1'b1;
    defparam \signature[164]~FF .SR_POLARITY = 1'b1;
    defparam \signature[164]~FF .D_POLARITY = 1'b1;
    defparam \signature[164]~FF .SR_SYNC = 1'b1;
    defparam \signature[164]~FF .SR_VALUE = 1'b0;
    defparam \signature[164]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[165]~FF  (.D(\useone/select_1071/Select_165/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[165] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[165]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[165]~FF .CE_POLARITY = 1'b1;
    defparam \signature[165]~FF .SR_POLARITY = 1'b1;
    defparam \signature[165]~FF .D_POLARITY = 1'b1;
    defparam \signature[165]~FF .SR_SYNC = 1'b1;
    defparam \signature[165]~FF .SR_VALUE = 1'b0;
    defparam \signature[165]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[166]~FF  (.D(\useone/select_1071/Select_166/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[166] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[166]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[166]~FF .CE_POLARITY = 1'b1;
    defparam \signature[166]~FF .SR_POLARITY = 1'b1;
    defparam \signature[166]~FF .D_POLARITY = 1'b1;
    defparam \signature[166]~FF .SR_SYNC = 1'b1;
    defparam \signature[166]~FF .SR_VALUE = 1'b0;
    defparam \signature[166]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[167]~FF  (.D(\useone/select_1071/Select_167/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[167] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[167]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[167]~FF .CE_POLARITY = 1'b1;
    defparam \signature[167]~FF .SR_POLARITY = 1'b1;
    defparam \signature[167]~FF .D_POLARITY = 1'b1;
    defparam \signature[167]~FF .SR_SYNC = 1'b1;
    defparam \signature[167]~FF .SR_VALUE = 1'b0;
    defparam \signature[167]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[168]~FF  (.D(\useone/select_1071/Select_168/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[168] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[168]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[168]~FF .CE_POLARITY = 1'b1;
    defparam \signature[168]~FF .SR_POLARITY = 1'b1;
    defparam \signature[168]~FF .D_POLARITY = 1'b1;
    defparam \signature[168]~FF .SR_SYNC = 1'b1;
    defparam \signature[168]~FF .SR_VALUE = 1'b0;
    defparam \signature[168]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[169]~FF  (.D(\useone/select_1071/Select_169/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[169] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[169]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[169]~FF .CE_POLARITY = 1'b1;
    defparam \signature[169]~FF .SR_POLARITY = 1'b1;
    defparam \signature[169]~FF .D_POLARITY = 1'b1;
    defparam \signature[169]~FF .SR_SYNC = 1'b1;
    defparam \signature[169]~FF .SR_VALUE = 1'b0;
    defparam \signature[169]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[170]~FF  (.D(\useone/select_1071/Select_170/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[170] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[170]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[170]~FF .CE_POLARITY = 1'b1;
    defparam \signature[170]~FF .SR_POLARITY = 1'b1;
    defparam \signature[170]~FF .D_POLARITY = 1'b1;
    defparam \signature[170]~FF .SR_SYNC = 1'b1;
    defparam \signature[170]~FF .SR_VALUE = 1'b0;
    defparam \signature[170]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[171]~FF  (.D(\useone/select_1071/Select_171/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[171] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[171]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[171]~FF .CE_POLARITY = 1'b1;
    defparam \signature[171]~FF .SR_POLARITY = 1'b1;
    defparam \signature[171]~FF .D_POLARITY = 1'b1;
    defparam \signature[171]~FF .SR_SYNC = 1'b1;
    defparam \signature[171]~FF .SR_VALUE = 1'b0;
    defparam \signature[171]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[172]~FF  (.D(\useone/select_1071/Select_172/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[172] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[172]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[172]~FF .CE_POLARITY = 1'b1;
    defparam \signature[172]~FF .SR_POLARITY = 1'b1;
    defparam \signature[172]~FF .D_POLARITY = 1'b1;
    defparam \signature[172]~FF .SR_SYNC = 1'b1;
    defparam \signature[172]~FF .SR_VALUE = 1'b0;
    defparam \signature[172]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[173]~FF  (.D(\useone/select_1071/Select_173/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[173] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[173]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[173]~FF .CE_POLARITY = 1'b1;
    defparam \signature[173]~FF .SR_POLARITY = 1'b1;
    defparam \signature[173]~FF .D_POLARITY = 1'b1;
    defparam \signature[173]~FF .SR_SYNC = 1'b1;
    defparam \signature[173]~FF .SR_VALUE = 1'b0;
    defparam \signature[173]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[174]~FF  (.D(\useone/select_1071/Select_174/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[174] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[174]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[174]~FF .CE_POLARITY = 1'b1;
    defparam \signature[174]~FF .SR_POLARITY = 1'b1;
    defparam \signature[174]~FF .D_POLARITY = 1'b1;
    defparam \signature[174]~FF .SR_SYNC = 1'b1;
    defparam \signature[174]~FF .SR_VALUE = 1'b0;
    defparam \signature[174]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[175]~FF  (.D(\useone/select_1071/Select_175/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[175] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[175]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[175]~FF .CE_POLARITY = 1'b1;
    defparam \signature[175]~FF .SR_POLARITY = 1'b1;
    defparam \signature[175]~FF .D_POLARITY = 1'b1;
    defparam \signature[175]~FF .SR_SYNC = 1'b1;
    defparam \signature[175]~FF .SR_VALUE = 1'b0;
    defparam \signature[175]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[176]~FF  (.D(\useone/select_1071/Select_176/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[176] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[176]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[176]~FF .CE_POLARITY = 1'b1;
    defparam \signature[176]~FF .SR_POLARITY = 1'b1;
    defparam \signature[176]~FF .D_POLARITY = 1'b1;
    defparam \signature[176]~FF .SR_SYNC = 1'b1;
    defparam \signature[176]~FF .SR_VALUE = 1'b0;
    defparam \signature[176]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[177]~FF  (.D(\useone/select_1071/Select_177/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[177] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[177]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[177]~FF .CE_POLARITY = 1'b1;
    defparam \signature[177]~FF .SR_POLARITY = 1'b1;
    defparam \signature[177]~FF .D_POLARITY = 1'b1;
    defparam \signature[177]~FF .SR_SYNC = 1'b1;
    defparam \signature[177]~FF .SR_VALUE = 1'b0;
    defparam \signature[177]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[178]~FF  (.D(\useone/select_1071/Select_178/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[178] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[178]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[178]~FF .CE_POLARITY = 1'b1;
    defparam \signature[178]~FF .SR_POLARITY = 1'b1;
    defparam \signature[178]~FF .D_POLARITY = 1'b1;
    defparam \signature[178]~FF .SR_SYNC = 1'b1;
    defparam \signature[178]~FF .SR_VALUE = 1'b0;
    defparam \signature[178]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[179]~FF  (.D(\useone/select_1071/Select_179/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[179] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[179]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[179]~FF .CE_POLARITY = 1'b1;
    defparam \signature[179]~FF .SR_POLARITY = 1'b1;
    defparam \signature[179]~FF .D_POLARITY = 1'b1;
    defparam \signature[179]~FF .SR_SYNC = 1'b1;
    defparam \signature[179]~FF .SR_VALUE = 1'b0;
    defparam \signature[179]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[180]~FF  (.D(\useone/select_1071/Select_180/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[180] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[180]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[180]~FF .CE_POLARITY = 1'b1;
    defparam \signature[180]~FF .SR_POLARITY = 1'b1;
    defparam \signature[180]~FF .D_POLARITY = 1'b1;
    defparam \signature[180]~FF .SR_SYNC = 1'b1;
    defparam \signature[180]~FF .SR_VALUE = 1'b0;
    defparam \signature[180]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[181]~FF  (.D(\useone/select_1071/Select_181/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[181] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[181]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[181]~FF .CE_POLARITY = 1'b1;
    defparam \signature[181]~FF .SR_POLARITY = 1'b1;
    defparam \signature[181]~FF .D_POLARITY = 1'b1;
    defparam \signature[181]~FF .SR_SYNC = 1'b1;
    defparam \signature[181]~FF .SR_VALUE = 1'b0;
    defparam \signature[181]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[182]~FF  (.D(\useone/select_1071/Select_182/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[182] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[182]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[182]~FF .CE_POLARITY = 1'b1;
    defparam \signature[182]~FF .SR_POLARITY = 1'b1;
    defparam \signature[182]~FF .D_POLARITY = 1'b1;
    defparam \signature[182]~FF .SR_SYNC = 1'b1;
    defparam \signature[182]~FF .SR_VALUE = 1'b0;
    defparam \signature[182]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[183]~FF  (.D(\useone/select_1071/Select_183/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[183] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[183]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[183]~FF .CE_POLARITY = 1'b1;
    defparam \signature[183]~FF .SR_POLARITY = 1'b1;
    defparam \signature[183]~FF .D_POLARITY = 1'b1;
    defparam \signature[183]~FF .SR_SYNC = 1'b1;
    defparam \signature[183]~FF .SR_VALUE = 1'b0;
    defparam \signature[183]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[184]~FF  (.D(\useone/select_1071/Select_184/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[184] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[184]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[184]~FF .CE_POLARITY = 1'b1;
    defparam \signature[184]~FF .SR_POLARITY = 1'b1;
    defparam \signature[184]~FF .D_POLARITY = 1'b1;
    defparam \signature[184]~FF .SR_SYNC = 1'b1;
    defparam \signature[184]~FF .SR_VALUE = 1'b0;
    defparam \signature[184]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[185]~FF  (.D(\useone/select_1071/Select_185/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[185] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[185]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[185]~FF .CE_POLARITY = 1'b1;
    defparam \signature[185]~FF .SR_POLARITY = 1'b1;
    defparam \signature[185]~FF .D_POLARITY = 1'b1;
    defparam \signature[185]~FF .SR_SYNC = 1'b1;
    defparam \signature[185]~FF .SR_VALUE = 1'b0;
    defparam \signature[185]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[186]~FF  (.D(\useone/select_1071/Select_186/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[186] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[186]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[186]~FF .CE_POLARITY = 1'b1;
    defparam \signature[186]~FF .SR_POLARITY = 1'b1;
    defparam \signature[186]~FF .D_POLARITY = 1'b1;
    defparam \signature[186]~FF .SR_SYNC = 1'b1;
    defparam \signature[186]~FF .SR_VALUE = 1'b0;
    defparam \signature[186]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[187]~FF  (.D(\useone/select_1071/Select_187/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[187] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[187]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[187]~FF .CE_POLARITY = 1'b1;
    defparam \signature[187]~FF .SR_POLARITY = 1'b1;
    defparam \signature[187]~FF .D_POLARITY = 1'b1;
    defparam \signature[187]~FF .SR_SYNC = 1'b1;
    defparam \signature[187]~FF .SR_VALUE = 1'b0;
    defparam \signature[187]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[188]~FF  (.D(\useone/select_1071/Select_188/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[188] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[188]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[188]~FF .CE_POLARITY = 1'b1;
    defparam \signature[188]~FF .SR_POLARITY = 1'b1;
    defparam \signature[188]~FF .D_POLARITY = 1'b1;
    defparam \signature[188]~FF .SR_SYNC = 1'b1;
    defparam \signature[188]~FF .SR_VALUE = 1'b0;
    defparam \signature[188]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[189]~FF  (.D(\useone/select_1071/Select_189/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[189] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[189]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[189]~FF .CE_POLARITY = 1'b1;
    defparam \signature[189]~FF .SR_POLARITY = 1'b1;
    defparam \signature[189]~FF .D_POLARITY = 1'b1;
    defparam \signature[189]~FF .SR_SYNC = 1'b1;
    defparam \signature[189]~FF .SR_VALUE = 1'b0;
    defparam \signature[189]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[190]~FF  (.D(\useone/select_1071/Select_190/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[190] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[190]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[190]~FF .CE_POLARITY = 1'b1;
    defparam \signature[190]~FF .SR_POLARITY = 1'b1;
    defparam \signature[190]~FF .D_POLARITY = 1'b1;
    defparam \signature[190]~FF .SR_SYNC = 1'b1;
    defparam \signature[190]~FF .SR_VALUE = 1'b0;
    defparam \signature[190]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[191]~FF  (.D(\useone/select_1071/Select_191/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[191] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[191]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[191]~FF .CE_POLARITY = 1'b1;
    defparam \signature[191]~FF .SR_POLARITY = 1'b1;
    defparam \signature[191]~FF .D_POLARITY = 1'b1;
    defparam \signature[191]~FF .SR_SYNC = 1'b1;
    defparam \signature[191]~FF .SR_VALUE = 1'b0;
    defparam \signature[191]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[192]~FF  (.D(\useone/select_1071/Select_192/n6 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[192] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[192]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[192]~FF .CE_POLARITY = 1'b1;
    defparam \signature[192]~FF .SR_POLARITY = 1'b1;
    defparam \signature[192]~FF .D_POLARITY = 1'b1;
    defparam \signature[192]~FF .SR_SYNC = 1'b1;
    defparam \signature[192]~FF .SR_VALUE = 1'b0;
    defparam \signature[192]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[193]~FF  (.D(\useone/select_1071/Select_193/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[193] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[193]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[193]~FF .CE_POLARITY = 1'b1;
    defparam \signature[193]~FF .SR_POLARITY = 1'b1;
    defparam \signature[193]~FF .D_POLARITY = 1'b1;
    defparam \signature[193]~FF .SR_SYNC = 1'b1;
    defparam \signature[193]~FF .SR_VALUE = 1'b0;
    defparam \signature[193]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[194]~FF  (.D(\useone/select_1071/Select_194/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[194] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[194]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[194]~FF .CE_POLARITY = 1'b1;
    defparam \signature[194]~FF .SR_POLARITY = 1'b1;
    defparam \signature[194]~FF .D_POLARITY = 1'b1;
    defparam \signature[194]~FF .SR_SYNC = 1'b1;
    defparam \signature[194]~FF .SR_VALUE = 1'b0;
    defparam \signature[194]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[195]~FF  (.D(\useone/select_1071/Select_195/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[195] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[195]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[195]~FF .CE_POLARITY = 1'b1;
    defparam \signature[195]~FF .SR_POLARITY = 1'b1;
    defparam \signature[195]~FF .D_POLARITY = 1'b1;
    defparam \signature[195]~FF .SR_SYNC = 1'b1;
    defparam \signature[195]~FF .SR_VALUE = 1'b0;
    defparam \signature[195]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[196]~FF  (.D(\useone/select_1071/Select_196/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[196] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[196]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[196]~FF .CE_POLARITY = 1'b1;
    defparam \signature[196]~FF .SR_POLARITY = 1'b1;
    defparam \signature[196]~FF .D_POLARITY = 1'b1;
    defparam \signature[196]~FF .SR_SYNC = 1'b1;
    defparam \signature[196]~FF .SR_VALUE = 1'b0;
    defparam \signature[196]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[197]~FF  (.D(\useone/select_1071/Select_197/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[197] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[197]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[197]~FF .CE_POLARITY = 1'b1;
    defparam \signature[197]~FF .SR_POLARITY = 1'b1;
    defparam \signature[197]~FF .D_POLARITY = 1'b1;
    defparam \signature[197]~FF .SR_SYNC = 1'b1;
    defparam \signature[197]~FF .SR_VALUE = 1'b0;
    defparam \signature[197]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[198]~FF  (.D(\useone/select_1071/Select_198/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[198] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[198]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[198]~FF .CE_POLARITY = 1'b1;
    defparam \signature[198]~FF .SR_POLARITY = 1'b1;
    defparam \signature[198]~FF .D_POLARITY = 1'b1;
    defparam \signature[198]~FF .SR_SYNC = 1'b1;
    defparam \signature[198]~FF .SR_VALUE = 1'b0;
    defparam \signature[198]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[199]~FF  (.D(\useone/select_1071/Select_199/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[199] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[199]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[199]~FF .CE_POLARITY = 1'b1;
    defparam \signature[199]~FF .SR_POLARITY = 1'b1;
    defparam \signature[199]~FF .D_POLARITY = 1'b1;
    defparam \signature[199]~FF .SR_SYNC = 1'b1;
    defparam \signature[199]~FF .SR_VALUE = 1'b0;
    defparam \signature[199]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[200]~FF  (.D(\useone/select_1071/Select_200/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[200] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[200]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[200]~FF .CE_POLARITY = 1'b1;
    defparam \signature[200]~FF .SR_POLARITY = 1'b1;
    defparam \signature[200]~FF .D_POLARITY = 1'b1;
    defparam \signature[200]~FF .SR_SYNC = 1'b1;
    defparam \signature[200]~FF .SR_VALUE = 1'b0;
    defparam \signature[200]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[201]~FF  (.D(\useone/select_1071/Select_201/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[201] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[201]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[201]~FF .CE_POLARITY = 1'b1;
    defparam \signature[201]~FF .SR_POLARITY = 1'b1;
    defparam \signature[201]~FF .D_POLARITY = 1'b1;
    defparam \signature[201]~FF .SR_SYNC = 1'b1;
    defparam \signature[201]~FF .SR_VALUE = 1'b0;
    defparam \signature[201]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[202]~FF  (.D(\useone/select_1071/Select_202/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[202] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[202]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[202]~FF .CE_POLARITY = 1'b1;
    defparam \signature[202]~FF .SR_POLARITY = 1'b1;
    defparam \signature[202]~FF .D_POLARITY = 1'b1;
    defparam \signature[202]~FF .SR_SYNC = 1'b1;
    defparam \signature[202]~FF .SR_VALUE = 1'b0;
    defparam \signature[202]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[203]~FF  (.D(\useone/select_1071/Select_203/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[203] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[203]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[203]~FF .CE_POLARITY = 1'b1;
    defparam \signature[203]~FF .SR_POLARITY = 1'b1;
    defparam \signature[203]~FF .D_POLARITY = 1'b1;
    defparam \signature[203]~FF .SR_SYNC = 1'b1;
    defparam \signature[203]~FF .SR_VALUE = 1'b0;
    defparam \signature[203]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[204]~FF  (.D(\useone/select_1071/Select_204/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[204] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[204]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[204]~FF .CE_POLARITY = 1'b1;
    defparam \signature[204]~FF .SR_POLARITY = 1'b1;
    defparam \signature[204]~FF .D_POLARITY = 1'b1;
    defparam \signature[204]~FF .SR_SYNC = 1'b1;
    defparam \signature[204]~FF .SR_VALUE = 1'b0;
    defparam \signature[204]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[205]~FF  (.D(\useone/select_1071/Select_205/n6 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[205] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[205]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[205]~FF .CE_POLARITY = 1'b1;
    defparam \signature[205]~FF .SR_POLARITY = 1'b1;
    defparam \signature[205]~FF .D_POLARITY = 1'b1;
    defparam \signature[205]~FF .SR_SYNC = 1'b1;
    defparam \signature[205]~FF .SR_VALUE = 1'b0;
    defparam \signature[205]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[206]~FF  (.D(\useone/select_1071/Select_206/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[206] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[206]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[206]~FF .CE_POLARITY = 1'b1;
    defparam \signature[206]~FF .SR_POLARITY = 1'b1;
    defparam \signature[206]~FF .D_POLARITY = 1'b1;
    defparam \signature[206]~FF .SR_SYNC = 1'b1;
    defparam \signature[206]~FF .SR_VALUE = 1'b0;
    defparam \signature[206]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[207]~FF  (.D(\useone/select_1071/Select_207/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[207] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[207]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[207]~FF .CE_POLARITY = 1'b1;
    defparam \signature[207]~FF .SR_POLARITY = 1'b1;
    defparam \signature[207]~FF .D_POLARITY = 1'b1;
    defparam \signature[207]~FF .SR_SYNC = 1'b1;
    defparam \signature[207]~FF .SR_VALUE = 1'b0;
    defparam \signature[207]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[208]~FF  (.D(\useone/select_1071/Select_208/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[208] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[208]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[208]~FF .CE_POLARITY = 1'b1;
    defparam \signature[208]~FF .SR_POLARITY = 1'b1;
    defparam \signature[208]~FF .D_POLARITY = 1'b1;
    defparam \signature[208]~FF .SR_SYNC = 1'b1;
    defparam \signature[208]~FF .SR_VALUE = 1'b0;
    defparam \signature[208]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[209]~FF  (.D(\useone/select_1071/Select_209/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[209] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[209]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[209]~FF .CE_POLARITY = 1'b1;
    defparam \signature[209]~FF .SR_POLARITY = 1'b1;
    defparam \signature[209]~FF .D_POLARITY = 1'b1;
    defparam \signature[209]~FF .SR_SYNC = 1'b1;
    defparam \signature[209]~FF .SR_VALUE = 1'b0;
    defparam \signature[209]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[210]~FF  (.D(\useone/select_1071/Select_210/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[210] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[210]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[210]~FF .CE_POLARITY = 1'b1;
    defparam \signature[210]~FF .SR_POLARITY = 1'b1;
    defparam \signature[210]~FF .D_POLARITY = 1'b1;
    defparam \signature[210]~FF .SR_SYNC = 1'b1;
    defparam \signature[210]~FF .SR_VALUE = 1'b0;
    defparam \signature[210]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[211]~FF  (.D(\useone/select_1071/Select_211/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[211] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[211]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[211]~FF .CE_POLARITY = 1'b1;
    defparam \signature[211]~FF .SR_POLARITY = 1'b1;
    defparam \signature[211]~FF .D_POLARITY = 1'b1;
    defparam \signature[211]~FF .SR_SYNC = 1'b1;
    defparam \signature[211]~FF .SR_VALUE = 1'b0;
    defparam \signature[211]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[212]~FF  (.D(\useone/select_1071/Select_212/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[212] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[212]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[212]~FF .CE_POLARITY = 1'b1;
    defparam \signature[212]~FF .SR_POLARITY = 1'b1;
    defparam \signature[212]~FF .D_POLARITY = 1'b1;
    defparam \signature[212]~FF .SR_SYNC = 1'b1;
    defparam \signature[212]~FF .SR_VALUE = 1'b0;
    defparam \signature[212]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[213]~FF  (.D(\useone/select_1071/Select_213/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[213] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[213]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[213]~FF .CE_POLARITY = 1'b1;
    defparam \signature[213]~FF .SR_POLARITY = 1'b1;
    defparam \signature[213]~FF .D_POLARITY = 1'b1;
    defparam \signature[213]~FF .SR_SYNC = 1'b1;
    defparam \signature[213]~FF .SR_VALUE = 1'b0;
    defparam \signature[213]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[214]~FF  (.D(\useone/select_1071/Select_214/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[214] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[214]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[214]~FF .CE_POLARITY = 1'b1;
    defparam \signature[214]~FF .SR_POLARITY = 1'b1;
    defparam \signature[214]~FF .D_POLARITY = 1'b1;
    defparam \signature[214]~FF .SR_SYNC = 1'b1;
    defparam \signature[214]~FF .SR_VALUE = 1'b0;
    defparam \signature[214]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[215]~FF  (.D(\useone/select_1071/Select_215/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[215] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[215]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[215]~FF .CE_POLARITY = 1'b1;
    defparam \signature[215]~FF .SR_POLARITY = 1'b1;
    defparam \signature[215]~FF .D_POLARITY = 1'b1;
    defparam \signature[215]~FF .SR_SYNC = 1'b1;
    defparam \signature[215]~FF .SR_VALUE = 1'b0;
    defparam \signature[215]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[216]~FF  (.D(\useone/select_1071/Select_216/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[216] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[216]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[216]~FF .CE_POLARITY = 1'b1;
    defparam \signature[216]~FF .SR_POLARITY = 1'b1;
    defparam \signature[216]~FF .D_POLARITY = 1'b1;
    defparam \signature[216]~FF .SR_SYNC = 1'b1;
    defparam \signature[216]~FF .SR_VALUE = 1'b0;
    defparam \signature[216]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[217]~FF  (.D(\useone/select_1071/Select_217/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[217] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[217]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[217]~FF .CE_POLARITY = 1'b1;
    defparam \signature[217]~FF .SR_POLARITY = 1'b1;
    defparam \signature[217]~FF .D_POLARITY = 1'b1;
    defparam \signature[217]~FF .SR_SYNC = 1'b1;
    defparam \signature[217]~FF .SR_VALUE = 1'b0;
    defparam \signature[217]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[218]~FF  (.D(\useone/select_1071/Select_218/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[218] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[218]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[218]~FF .CE_POLARITY = 1'b1;
    defparam \signature[218]~FF .SR_POLARITY = 1'b1;
    defparam \signature[218]~FF .D_POLARITY = 1'b1;
    defparam \signature[218]~FF .SR_SYNC = 1'b1;
    defparam \signature[218]~FF .SR_VALUE = 1'b0;
    defparam \signature[218]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[219]~FF  (.D(\useone/select_1071/Select_219/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[219] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[219]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[219]~FF .CE_POLARITY = 1'b1;
    defparam \signature[219]~FF .SR_POLARITY = 1'b1;
    defparam \signature[219]~FF .D_POLARITY = 1'b1;
    defparam \signature[219]~FF .SR_SYNC = 1'b1;
    defparam \signature[219]~FF .SR_VALUE = 1'b0;
    defparam \signature[219]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[220]~FF  (.D(\useone/select_1071/Select_220/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[220] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[220]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[220]~FF .CE_POLARITY = 1'b1;
    defparam \signature[220]~FF .SR_POLARITY = 1'b1;
    defparam \signature[220]~FF .D_POLARITY = 1'b1;
    defparam \signature[220]~FF .SR_SYNC = 1'b1;
    defparam \signature[220]~FF .SR_VALUE = 1'b0;
    defparam \signature[220]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[221]~FF  (.D(\useone/select_1071/Select_221/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[221] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[221]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[221]~FF .CE_POLARITY = 1'b1;
    defparam \signature[221]~FF .SR_POLARITY = 1'b1;
    defparam \signature[221]~FF .D_POLARITY = 1'b1;
    defparam \signature[221]~FF .SR_SYNC = 1'b1;
    defparam \signature[221]~FF .SR_VALUE = 1'b0;
    defparam \signature[221]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[222]~FF  (.D(\useone/select_1071/Select_222/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[222] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[222]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[222]~FF .CE_POLARITY = 1'b1;
    defparam \signature[222]~FF .SR_POLARITY = 1'b1;
    defparam \signature[222]~FF .D_POLARITY = 1'b1;
    defparam \signature[222]~FF .SR_SYNC = 1'b1;
    defparam \signature[222]~FF .SR_VALUE = 1'b0;
    defparam \signature[222]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[223]~FF  (.D(\useone/select_1071/Select_223/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[223] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[223]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[223]~FF .CE_POLARITY = 1'b1;
    defparam \signature[223]~FF .SR_POLARITY = 1'b1;
    defparam \signature[223]~FF .D_POLARITY = 1'b1;
    defparam \signature[223]~FF .SR_SYNC = 1'b1;
    defparam \signature[223]~FF .SR_VALUE = 1'b0;
    defparam \signature[223]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[224]~FF  (.D(\useone/select_1071/Select_224/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[224] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[224]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[224]~FF .CE_POLARITY = 1'b1;
    defparam \signature[224]~FF .SR_POLARITY = 1'b1;
    defparam \signature[224]~FF .D_POLARITY = 1'b1;
    defparam \signature[224]~FF .SR_SYNC = 1'b1;
    defparam \signature[224]~FF .SR_VALUE = 1'b0;
    defparam \signature[224]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[225]~FF  (.D(\useone/select_1071/Select_225/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[225] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[225]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[225]~FF .CE_POLARITY = 1'b1;
    defparam \signature[225]~FF .SR_POLARITY = 1'b1;
    defparam \signature[225]~FF .D_POLARITY = 1'b1;
    defparam \signature[225]~FF .SR_SYNC = 1'b1;
    defparam \signature[225]~FF .SR_VALUE = 1'b0;
    defparam \signature[225]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[226]~FF  (.D(\useone/select_1071/Select_226/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[226] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[226]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[226]~FF .CE_POLARITY = 1'b1;
    defparam \signature[226]~FF .SR_POLARITY = 1'b1;
    defparam \signature[226]~FF .D_POLARITY = 1'b1;
    defparam \signature[226]~FF .SR_SYNC = 1'b1;
    defparam \signature[226]~FF .SR_VALUE = 1'b0;
    defparam \signature[226]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[227]~FF  (.D(\useone/select_1071/Select_227/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[227] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[227]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[227]~FF .CE_POLARITY = 1'b1;
    defparam \signature[227]~FF .SR_POLARITY = 1'b1;
    defparam \signature[227]~FF .D_POLARITY = 1'b1;
    defparam \signature[227]~FF .SR_SYNC = 1'b1;
    defparam \signature[227]~FF .SR_VALUE = 1'b0;
    defparam \signature[227]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[228]~FF  (.D(\useone/select_1071/Select_228/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[228] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[228]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[228]~FF .CE_POLARITY = 1'b1;
    defparam \signature[228]~FF .SR_POLARITY = 1'b1;
    defparam \signature[228]~FF .D_POLARITY = 1'b1;
    defparam \signature[228]~FF .SR_SYNC = 1'b1;
    defparam \signature[228]~FF .SR_VALUE = 1'b0;
    defparam \signature[228]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[229]~FF  (.D(\useone/select_1071/Select_229/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[229] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[229]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[229]~FF .CE_POLARITY = 1'b1;
    defparam \signature[229]~FF .SR_POLARITY = 1'b1;
    defparam \signature[229]~FF .D_POLARITY = 1'b1;
    defparam \signature[229]~FF .SR_SYNC = 1'b1;
    defparam \signature[229]~FF .SR_VALUE = 1'b0;
    defparam \signature[229]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[230]~FF  (.D(\useone/select_1071/Select_230/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[230] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[230]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[230]~FF .CE_POLARITY = 1'b1;
    defparam \signature[230]~FF .SR_POLARITY = 1'b1;
    defparam \signature[230]~FF .D_POLARITY = 1'b1;
    defparam \signature[230]~FF .SR_SYNC = 1'b1;
    defparam \signature[230]~FF .SR_VALUE = 1'b0;
    defparam \signature[230]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[231]~FF  (.D(\useone/select_1071/Select_231/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[231] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[231]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[231]~FF .CE_POLARITY = 1'b1;
    defparam \signature[231]~FF .SR_POLARITY = 1'b1;
    defparam \signature[231]~FF .D_POLARITY = 1'b1;
    defparam \signature[231]~FF .SR_SYNC = 1'b1;
    defparam \signature[231]~FF .SR_VALUE = 1'b0;
    defparam \signature[231]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[232]~FF  (.D(\useone/select_1071/Select_232/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[232] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[232]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[232]~FF .CE_POLARITY = 1'b1;
    defparam \signature[232]~FF .SR_POLARITY = 1'b1;
    defparam \signature[232]~FF .D_POLARITY = 1'b1;
    defparam \signature[232]~FF .SR_SYNC = 1'b1;
    defparam \signature[232]~FF .SR_VALUE = 1'b0;
    defparam \signature[232]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[233]~FF  (.D(\useone/select_1071/Select_233/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[233] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[233]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[233]~FF .CE_POLARITY = 1'b1;
    defparam \signature[233]~FF .SR_POLARITY = 1'b1;
    defparam \signature[233]~FF .D_POLARITY = 1'b1;
    defparam \signature[233]~FF .SR_SYNC = 1'b1;
    defparam \signature[233]~FF .SR_VALUE = 1'b0;
    defparam \signature[233]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[234]~FF  (.D(\useone/select_1071/Select_234/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[234] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[234]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[234]~FF .CE_POLARITY = 1'b1;
    defparam \signature[234]~FF .SR_POLARITY = 1'b1;
    defparam \signature[234]~FF .D_POLARITY = 1'b1;
    defparam \signature[234]~FF .SR_SYNC = 1'b1;
    defparam \signature[234]~FF .SR_VALUE = 1'b0;
    defparam \signature[234]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[235]~FF  (.D(\useone/select_1071/Select_235/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[235] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[235]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[235]~FF .CE_POLARITY = 1'b1;
    defparam \signature[235]~FF .SR_POLARITY = 1'b1;
    defparam \signature[235]~FF .D_POLARITY = 1'b1;
    defparam \signature[235]~FF .SR_SYNC = 1'b1;
    defparam \signature[235]~FF .SR_VALUE = 1'b0;
    defparam \signature[235]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[236]~FF  (.D(\useone/select_1071/Select_236/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[236] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[236]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[236]~FF .CE_POLARITY = 1'b1;
    defparam \signature[236]~FF .SR_POLARITY = 1'b1;
    defparam \signature[236]~FF .D_POLARITY = 1'b1;
    defparam \signature[236]~FF .SR_SYNC = 1'b1;
    defparam \signature[236]~FF .SR_VALUE = 1'b0;
    defparam \signature[236]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[237]~FF  (.D(\useone/select_1071/Select_237/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[237] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[237]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[237]~FF .CE_POLARITY = 1'b1;
    defparam \signature[237]~FF .SR_POLARITY = 1'b1;
    defparam \signature[237]~FF .D_POLARITY = 1'b1;
    defparam \signature[237]~FF .SR_SYNC = 1'b1;
    defparam \signature[237]~FF .SR_VALUE = 1'b0;
    defparam \signature[237]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[238]~FF  (.D(\useone/select_1071/Select_238/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[238] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[238]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[238]~FF .CE_POLARITY = 1'b1;
    defparam \signature[238]~FF .SR_POLARITY = 1'b1;
    defparam \signature[238]~FF .D_POLARITY = 1'b1;
    defparam \signature[238]~FF .SR_SYNC = 1'b1;
    defparam \signature[238]~FF .SR_VALUE = 1'b0;
    defparam \signature[238]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[239]~FF  (.D(\useone/select_1071/Select_239/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[239] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[239]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[239]~FF .CE_POLARITY = 1'b1;
    defparam \signature[239]~FF .SR_POLARITY = 1'b1;
    defparam \signature[239]~FF .D_POLARITY = 1'b1;
    defparam \signature[239]~FF .SR_SYNC = 1'b1;
    defparam \signature[239]~FF .SR_VALUE = 1'b0;
    defparam \signature[239]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[240]~FF  (.D(\useone/select_1071/Select_240/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[240] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[240]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[240]~FF .CE_POLARITY = 1'b1;
    defparam \signature[240]~FF .SR_POLARITY = 1'b1;
    defparam \signature[240]~FF .D_POLARITY = 1'b1;
    defparam \signature[240]~FF .SR_SYNC = 1'b1;
    defparam \signature[240]~FF .SR_VALUE = 1'b0;
    defparam \signature[240]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[241]~FF  (.D(\useone/select_1071/Select_241/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[241] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[241]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[241]~FF .CE_POLARITY = 1'b1;
    defparam \signature[241]~FF .SR_POLARITY = 1'b1;
    defparam \signature[241]~FF .D_POLARITY = 1'b1;
    defparam \signature[241]~FF .SR_SYNC = 1'b1;
    defparam \signature[241]~FF .SR_VALUE = 1'b0;
    defparam \signature[241]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[242]~FF  (.D(\useone/select_1071/Select_242/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[242] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[242]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[242]~FF .CE_POLARITY = 1'b1;
    defparam \signature[242]~FF .SR_POLARITY = 1'b1;
    defparam \signature[242]~FF .D_POLARITY = 1'b1;
    defparam \signature[242]~FF .SR_SYNC = 1'b1;
    defparam \signature[242]~FF .SR_VALUE = 1'b0;
    defparam \signature[242]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[243]~FF  (.D(\useone/select_1071/Select_243/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[243] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[243]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[243]~FF .CE_POLARITY = 1'b1;
    defparam \signature[243]~FF .SR_POLARITY = 1'b1;
    defparam \signature[243]~FF .D_POLARITY = 1'b1;
    defparam \signature[243]~FF .SR_SYNC = 1'b1;
    defparam \signature[243]~FF .SR_VALUE = 1'b0;
    defparam \signature[243]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[244]~FF  (.D(\useone/select_1071/Select_244/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[244] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[244]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[244]~FF .CE_POLARITY = 1'b1;
    defparam \signature[244]~FF .SR_POLARITY = 1'b1;
    defparam \signature[244]~FF .D_POLARITY = 1'b1;
    defparam \signature[244]~FF .SR_SYNC = 1'b1;
    defparam \signature[244]~FF .SR_VALUE = 1'b0;
    defparam \signature[244]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[245]~FF  (.D(\useone/select_1071/Select_245/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[245] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[245]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[245]~FF .CE_POLARITY = 1'b1;
    defparam \signature[245]~FF .SR_POLARITY = 1'b1;
    defparam \signature[245]~FF .D_POLARITY = 1'b1;
    defparam \signature[245]~FF .SR_SYNC = 1'b1;
    defparam \signature[245]~FF .SR_VALUE = 1'b0;
    defparam \signature[245]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[246]~FF  (.D(\useone/select_1071/Select_246/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[246] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[246]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[246]~FF .CE_POLARITY = 1'b1;
    defparam \signature[246]~FF .SR_POLARITY = 1'b1;
    defparam \signature[246]~FF .D_POLARITY = 1'b1;
    defparam \signature[246]~FF .SR_SYNC = 1'b1;
    defparam \signature[246]~FF .SR_VALUE = 1'b0;
    defparam \signature[246]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[247]~FF  (.D(\useone/select_1071/Select_247/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[247] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[247]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[247]~FF .CE_POLARITY = 1'b1;
    defparam \signature[247]~FF .SR_POLARITY = 1'b1;
    defparam \signature[247]~FF .D_POLARITY = 1'b1;
    defparam \signature[247]~FF .SR_SYNC = 1'b1;
    defparam \signature[247]~FF .SR_VALUE = 1'b0;
    defparam \signature[247]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[248]~FF  (.D(\useone/select_1071/Select_248/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[248] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[248]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[248]~FF .CE_POLARITY = 1'b1;
    defparam \signature[248]~FF .SR_POLARITY = 1'b1;
    defparam \signature[248]~FF .D_POLARITY = 1'b1;
    defparam \signature[248]~FF .SR_SYNC = 1'b1;
    defparam \signature[248]~FF .SR_VALUE = 1'b0;
    defparam \signature[248]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[249]~FF  (.D(\useone/select_1071/Select_249/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[249] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[249]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[249]~FF .CE_POLARITY = 1'b1;
    defparam \signature[249]~FF .SR_POLARITY = 1'b1;
    defparam \signature[249]~FF .D_POLARITY = 1'b1;
    defparam \signature[249]~FF .SR_SYNC = 1'b1;
    defparam \signature[249]~FF .SR_VALUE = 1'b0;
    defparam \signature[249]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[250]~FF  (.D(\useone/select_1071/Select_250/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[250] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[250]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[250]~FF .CE_POLARITY = 1'b1;
    defparam \signature[250]~FF .SR_POLARITY = 1'b1;
    defparam \signature[250]~FF .D_POLARITY = 1'b1;
    defparam \signature[250]~FF .SR_SYNC = 1'b1;
    defparam \signature[250]~FF .SR_VALUE = 1'b0;
    defparam \signature[250]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[251]~FF  (.D(\useone/select_1071/Select_251/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[251] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[251]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[251]~FF .CE_POLARITY = 1'b1;
    defparam \signature[251]~FF .SR_POLARITY = 1'b1;
    defparam \signature[251]~FF .D_POLARITY = 1'b1;
    defparam \signature[251]~FF .SR_SYNC = 1'b1;
    defparam \signature[251]~FF .SR_VALUE = 1'b0;
    defparam \signature[251]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[252]~FF  (.D(\useone/select_1071/Select_252/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[252] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[252]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[252]~FF .CE_POLARITY = 1'b1;
    defparam \signature[252]~FF .SR_POLARITY = 1'b1;
    defparam \signature[252]~FF .D_POLARITY = 1'b1;
    defparam \signature[252]~FF .SR_SYNC = 1'b1;
    defparam \signature[252]~FF .SR_VALUE = 1'b0;
    defparam \signature[252]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[253]~FF  (.D(\useone/select_1071/Select_253/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[253] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[253]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[253]~FF .CE_POLARITY = 1'b1;
    defparam \signature[253]~FF .SR_POLARITY = 1'b1;
    defparam \signature[253]~FF .D_POLARITY = 1'b1;
    defparam \signature[253]~FF .SR_SYNC = 1'b1;
    defparam \signature[253]~FF .SR_VALUE = 1'b0;
    defparam \signature[253]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[254]~FF  (.D(\useone/select_1071/Select_254/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[254] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[254]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[254]~FF .CE_POLARITY = 1'b1;
    defparam \signature[254]~FF .SR_POLARITY = 1'b1;
    defparam \signature[254]~FF .D_POLARITY = 1'b1;
    defparam \signature[254]~FF .SR_SYNC = 1'b1;
    defparam \signature[254]~FF .SR_VALUE = 1'b0;
    defparam \signature[254]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \signature[255]~FF  (.D(\useone/select_1071/Select_255/n2 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\signature[255] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(240)
    defparam \signature[255]~FF .CLK_POLARITY = 1'b1;
    defparam \signature[255]~FF .CE_POLARITY = 1'b1;
    defparam \signature[255]~FF .SR_POLARITY = 1'b1;
    defparam \signature[255]~FF .D_POLARITY = 1'b1;
    defparam \signature[255]~FF .SR_SYNC = 1'b1;
    defparam \signature[255]~FF .SR_VALUE = 1'b0;
    defparam \signature[255]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[0]~FF  (.D(\useuart/n844 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[0]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[0]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[0]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[0]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[0]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_uart_tx_2~FF  (.D(\useuart/n634 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(o_uart_tx_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \o_uart_tx_2~FF .CLK_POLARITY = 1'b1;
    defparam \o_uart_tx_2~FF .CE_POLARITY = 1'b0;
    defparam \o_uart_tx_2~FF .SR_POLARITY = 1'b1;
    defparam \o_uart_tx_2~FF .D_POLARITY = 1'b0;
    defparam \o_uart_tx_2~FF .SR_SYNC = 1'b1;
    defparam \o_uart_tx_2~FF .SR_VALUE = 1'b0;
    defparam \o_uart_tx_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Bit_Index[0]~FF  (.D(\useuart/n848 ), .CE(ceg_net79), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Bit_Index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Bit_Index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[0]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Bit_Index[0]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[0]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[0]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Bit_Index[0]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Bit_Index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \o_Tx_active~FF  (.D(\useuart/r_SM_Main[1] ), .CE(ceg_net77), 
           .CLK(\clk~O ), .SR(1'b0), .Q(o_Tx_active)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \o_Tx_active~FF .CLK_POLARITY = 1'b1;
    defparam \o_Tx_active~FF .CE_POLARITY = 1'b0;
    defparam \o_Tx_active~FF .SR_POLARITY = 1'b1;
    defparam \o_Tx_active~FF .D_POLARITY = 1'b0;
    defparam \o_Tx_active~FF .SR_SYNC = 1'b1;
    defparam \o_Tx_active~FF .SR_VALUE = 1'b0;
    defparam \o_Tx_active~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Tx_Data[0]~FF  (.D(\data_chunk[0] ), .CE(\useuart/n960 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Tx_Data[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Tx_Data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[0]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[0]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[0]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[0]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Tx_Data[0]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Tx_Data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_SM_Main[0]~FF  (.D(\useuart/n840 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\useuart/r_SM_Main[2] ), .Q(\useuart/r_SM_Main[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_SM_Main[0]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[0]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[0]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[0]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[0]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_SM_Main[0]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_SM_Main[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[1]~FF  (.D(\useuart/n708 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[1]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[1]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[1]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[1]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[1]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[2]~FF  (.D(\useuart/n711 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[2]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[2]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[2]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[2]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[2]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[3]~FF  (.D(\useuart/n714 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[3]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[3]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[3]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[3]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[3]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[4]~FF  (.D(\useuart/n717 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[4]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[4]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[4]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[4]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[4]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[5]~FF  (.D(\useuart/n720 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[5]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[5]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[5]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[5]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[5]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[6]~FF  (.D(\useuart/n723 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[6]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[6]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[6]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[6]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[6]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[7]~FF  (.D(\useuart/n726 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[7]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[7]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[7]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[7]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[7]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[8]~FF  (.D(\useuart/n729 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[8]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[8]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[8]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[8]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[8]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[8]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[9]~FF  (.D(\useuart/n732 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[9]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[9]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[9]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[9]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[9]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[9]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[10]~FF  (.D(\useuart/n735 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[10]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[10]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[10]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[10]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[10]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[10]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[11]~FF  (.D(\useuart/n738 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[11]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[11]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[11]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[11]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[11]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[11]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Clock_Count[12]~FF  (.D(\useuart/n741 ), .CE(\useuart/r_SM_Main[2] ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Clock_Count[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Clock_Count[12]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[12]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Clock_Count[12]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[12]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Clock_Count[12]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Clock_Count[12]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Clock_Count[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Bit_Index[1]~FF  (.D(\useuart/n802 ), .CE(ceg_net79), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Bit_Index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Bit_Index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[1]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Bit_Index[1]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[1]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[1]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Bit_Index[1]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Bit_Index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Bit_Index[2]~FF  (.D(\useuart/n806 ), .CE(ceg_net79), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Bit_Index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Bit_Index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[2]~FF .CE_POLARITY = 1'b0;
    defparam \useuart/r_Bit_Index[2]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[2]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Bit_Index[2]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Bit_Index[2]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Bit_Index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Tx_Data[1]~FF  (.D(\data_chunk[1] ), .CE(\useuart/n960 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Tx_Data[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Tx_Data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[1]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[1]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[1]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[1]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Tx_Data[1]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Tx_Data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Tx_Data[2]~FF  (.D(\data_chunk[2] ), .CE(\useuart/n960 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Tx_Data[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Tx_Data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[2]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[2]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[2]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[2]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Tx_Data[2]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Tx_Data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Tx_Data[3]~FF  (.D(\data_chunk[3] ), .CE(\useuart/n960 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Tx_Data[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Tx_Data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[3]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[3]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[3]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[3]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Tx_Data[3]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Tx_Data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Tx_Data[4]~FF  (.D(\data_chunk[4] ), .CE(\useuart/n960 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Tx_Data[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Tx_Data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[4]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[4]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[4]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[4]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Tx_Data[4]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Tx_Data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Tx_Data[5]~FF  (.D(\data_chunk[5] ), .CE(\useuart/n960 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Tx_Data[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Tx_Data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[5]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[5]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[5]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[5]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Tx_Data[5]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Tx_Data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Tx_Data[6]~FF  (.D(\data_chunk[6] ), .CE(\useuart/n960 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Tx_Data[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Tx_Data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[6]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[6]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[6]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[6]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Tx_Data[6]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Tx_Data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_Tx_Data[7]~FF  (.D(\data_chunk[7] ), .CE(\useuart/n960 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\useuart/r_Tx_Data[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_Tx_Data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[7]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[7]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[7]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_Tx_Data[7]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_Tx_Data[7]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_Tx_Data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_SM_Main[1]~FF  (.D(\useuart/n836 ), .CE(1'b1), .CLK(\clk~O ), 
           .SR(\useuart/r_SM_Main[2] ), .Q(\useuart/r_SM_Main[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_SM_Main[1]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[1]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[1]~FF .SR_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[1]~FF .D_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[1]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_SM_Main[1]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_SM_Main[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \useuart/r_SM_Main[2]~FF  (.D(\useuart/LessThan_9/n26 ), .CE(1'b1), 
           .CLK(\clk~O ), .SR(\useuart/n942 ), .Q(\useuart/r_SM_Main[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\uart_tx.sv(114)
    defparam \useuart/r_SM_Main[2]~FF .CLK_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[2]~FF .CE_POLARITY = 1'b1;
    defparam \useuart/r_SM_Main[2]~FF .SR_POLARITY = 1'b0;
    defparam \useuart/r_SM_Main[2]~FF .D_POLARITY = 1'b0;
    defparam \useuart/r_SM_Main[2]~FF .SR_SYNC = 1'b1;
    defparam \useuart/r_SM_Main[2]~FF .SR_VALUE = 1'b0;
    defparam \useuart/r_SM_Main[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \chunk_index[1]~FF  (.D(n935_2), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\chunk_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \chunk_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \chunk_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \chunk_index[1]~FF .SR_POLARITY = 1'b1;
    defparam \chunk_index[1]~FF .D_POLARITY = 1'b1;
    defparam \chunk_index[1]~FF .SR_SYNC = 1'b0;
    defparam \chunk_index[1]~FF .SR_VALUE = 1'b0;
    defparam \chunk_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \chunk_index[2]~FF  (.D(n940_2), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\chunk_index[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \chunk_index[2]~FF .CLK_POLARITY = 1'b1;
    defparam \chunk_index[2]~FF .CE_POLARITY = 1'b0;
    defparam \chunk_index[2]~FF .SR_POLARITY = 1'b1;
    defparam \chunk_index[2]~FF .D_POLARITY = 1'b1;
    defparam \chunk_index[2]~FF .SR_SYNC = 1'b0;
    defparam \chunk_index[2]~FF .SR_VALUE = 1'b0;
    defparam \chunk_index[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \chunk_index[3]~FF  (.D(n945_2), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\chunk_index[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \chunk_index[3]~FF .CLK_POLARITY = 1'b1;
    defparam \chunk_index[3]~FF .CE_POLARITY = 1'b0;
    defparam \chunk_index[3]~FF .SR_POLARITY = 1'b1;
    defparam \chunk_index[3]~FF .D_POLARITY = 1'b1;
    defparam \chunk_index[3]~FF .SR_SYNC = 1'b0;
    defparam \chunk_index[3]~FF .SR_VALUE = 1'b0;
    defparam \chunk_index[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \chunk_index[4]~FF  (.D(n950_2), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\chunk_index[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \chunk_index[4]~FF .CLK_POLARITY = 1'b1;
    defparam \chunk_index[4]~FF .CE_POLARITY = 1'b0;
    defparam \chunk_index[4]~FF .SR_POLARITY = 1'b1;
    defparam \chunk_index[4]~FF .D_POLARITY = 1'b1;
    defparam \chunk_index[4]~FF .SR_SYNC = 1'b0;
    defparam \chunk_index[4]~FF .SR_VALUE = 1'b0;
    defparam \chunk_index[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \chunk_index[5]~FF  (.D(n955_2), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\chunk_index[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \chunk_index[5]~FF .CLK_POLARITY = 1'b1;
    defparam \chunk_index[5]~FF .CE_POLARITY = 1'b0;
    defparam \chunk_index[5]~FF .SR_POLARITY = 1'b1;
    defparam \chunk_index[5]~FF .D_POLARITY = 1'b1;
    defparam \chunk_index[5]~FF .SR_SYNC = 1'b0;
    defparam \chunk_index[5]~FF .SR_VALUE = 1'b0;
    defparam \chunk_index[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \state[1]~FF  (.D(n868_2), .CE(ceg_net99), .CLK(\clk~O ), .SR(rst), 
           .Q(\state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \state[1]~FF .CE_POLARITY = 1'b0;
    defparam \state[1]~FF .SR_POLARITY = 1'b1;
    defparam \state[1]~FF .D_POLARITY = 1'b1;
    defparam \state[1]~FF .SR_SYNC = 1'b0;
    defparam \state[1]~FF .SR_VALUE = 1'b0;
    defparam \state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_chunk[1]~FF  (.D(n827), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\data_chunk[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \data_chunk[1]~FF .CLK_POLARITY = 1'b1;
    defparam \data_chunk[1]~FF .CE_POLARITY = 1'b0;
    defparam \data_chunk[1]~FF .SR_POLARITY = 1'b1;
    defparam \data_chunk[1]~FF .D_POLARITY = 1'b1;
    defparam \data_chunk[1]~FF .SR_SYNC = 1'b0;
    defparam \data_chunk[1]~FF .SR_VALUE = 1'b0;
    defparam \data_chunk[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_chunk[2]~FF  (.D(n826), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\data_chunk[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \data_chunk[2]~FF .CLK_POLARITY = 1'b1;
    defparam \data_chunk[2]~FF .CE_POLARITY = 1'b0;
    defparam \data_chunk[2]~FF .SR_POLARITY = 1'b1;
    defparam \data_chunk[2]~FF .D_POLARITY = 1'b1;
    defparam \data_chunk[2]~FF .SR_SYNC = 1'b0;
    defparam \data_chunk[2]~FF .SR_VALUE = 1'b0;
    defparam \data_chunk[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_chunk[3]~FF  (.D(n825), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\data_chunk[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \data_chunk[3]~FF .CLK_POLARITY = 1'b1;
    defparam \data_chunk[3]~FF .CE_POLARITY = 1'b0;
    defparam \data_chunk[3]~FF .SR_POLARITY = 1'b1;
    defparam \data_chunk[3]~FF .D_POLARITY = 1'b1;
    defparam \data_chunk[3]~FF .SR_SYNC = 1'b0;
    defparam \data_chunk[3]~FF .SR_VALUE = 1'b0;
    defparam \data_chunk[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_chunk[4]~FF  (.D(n824), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\data_chunk[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \data_chunk[4]~FF .CLK_POLARITY = 1'b1;
    defparam \data_chunk[4]~FF .CE_POLARITY = 1'b0;
    defparam \data_chunk[4]~FF .SR_POLARITY = 1'b1;
    defparam \data_chunk[4]~FF .D_POLARITY = 1'b1;
    defparam \data_chunk[4]~FF .SR_SYNC = 1'b0;
    defparam \data_chunk[4]~FF .SR_VALUE = 1'b0;
    defparam \data_chunk[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_chunk[5]~FF  (.D(n823), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\data_chunk[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \data_chunk[5]~FF .CLK_POLARITY = 1'b1;
    defparam \data_chunk[5]~FF .CE_POLARITY = 1'b0;
    defparam \data_chunk[5]~FF .SR_POLARITY = 1'b1;
    defparam \data_chunk[5]~FF .D_POLARITY = 1'b1;
    defparam \data_chunk[5]~FF .SR_SYNC = 1'b0;
    defparam \data_chunk[5]~FF .SR_VALUE = 1'b0;
    defparam \data_chunk[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_chunk[6]~FF  (.D(n822), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\data_chunk[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \data_chunk[6]~FF .CLK_POLARITY = 1'b1;
    defparam \data_chunk[6]~FF .CE_POLARITY = 1'b0;
    defparam \data_chunk[6]~FF .SR_POLARITY = 1'b1;
    defparam \data_chunk[6]~FF .D_POLARITY = 1'b1;
    defparam \data_chunk[6]~FF .SR_SYNC = 1'b0;
    defparam \data_chunk[6]~FF .SR_VALUE = 1'b0;
    defparam \data_chunk[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \data_chunk[7]~FF  (.D(n821), .CE(ceg_net40), .CLK(\clk~O ), 
           .SR(rst), .Q(\data_chunk[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\top.sv(83)
    defparam \data_chunk[7]~FF .CLK_POLARITY = 1'b1;
    defparam \data_chunk[7]~FF .CE_POLARITY = 1'b0;
    defparam \data_chunk[7]~FF .SR_POLARITY = 1'b1;
    defparam \data_chunk[7]~FF .D_POLARITY = 1'b1;
    defparam \data_chunk[7]~FF .SR_SYNC = 1'b0;
    defparam \data_chunk[7]~FF .SR_VALUE = 1'b0;
    defparam \data_chunk[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \i131/useone/w[17][23]~FF  (.D(n1191_2), .CE(\useone/equal_1067/n7 ), 
           .CLK(\clk~O ), .SR(1'b0), .Q(\i131/useone/w[17][23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(18)
    defparam \i131/useone/w[17][23]~FF .CLK_POLARITY = 1'b1;
    defparam \i131/useone/w[17][23]~FF .CE_POLARITY = 1'b0;
    defparam \i131/useone/w[17][23]~FF .SR_POLARITY = 1'b1;
    defparam \i131/useone/w[17][23]~FF .D_POLARITY = 1'b1;
    defparam \i131/useone/w[17][23]~FF .SR_SYNC = 1'b1;
    defparam \i131/useone/w[17][23]~FF .SR_VALUE = 1'b0;
    defparam \i131/useone/w[17][23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \useone/add_995/i1  (.I0(\useone/h[0] ), .I1(n1790), .CI(1'b0), 
            .O(n10), .CO(n11)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i1 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i1  (.I0(n10), .I1(n1792), .CI(1'b0), .O(n12), 
            .CO(n13)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i1  (.I0(n12), .I1(n1794), .CI(1'b0), .O(n14), 
            .CO(n15)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i1  (.I0(n14), .I1(n1796), .CI(1'b0), .O(n16), 
            .CO(n17)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i1  (.I0(n1797), .I1(n1798), .CI(1'b0), .O(n18), 
            .CO(n19)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i1  (.I0(\useone/d[0] ), .I1(n16), .CI(1'b0), 
            .O(n20), .CO(n21)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i1  (.I0(n16), .I1(n18), .CI(1'b0), .O(n22), 
            .CO(n23)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i1  (.I0(\useone/H0[0] ), .I1(\useone/a[0] ), 
            .CI(1'b0), .O(n24), .CO(n25)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i1 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i1  (.I0(\useone/H1[0] ), .I1(\useone/b[0] ), 
            .CI(1'b0), .O(n26), .CO(n27)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i1 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i1  (.I0(\useone/H2[0] ), .I1(\useone/c[0] ), 
            .CI(1'b0), .O(n28), .CO(n29)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i1  (.I0(\useone/H3[0] ), .I1(\useone/d[0] ), 
            .CI(1'b0), .O(n30), .CO(n31)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i1  (.I0(\useone/H4[0] ), .I1(\useone/e[0] ), 
            .CI(1'b0), .O(n32), .CO(n33)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i1 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i1  (.I0(\useone/H5[0] ), .I1(\useone/f[0] ), 
            .CI(1'b0), .O(n34), .CO(n35)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i1 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i1  (.I0(\useone/H6[0] ), .I1(\useone/g[0] ), 
            .CI(1'b0), .O(n36), .CO(n37)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i1 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i1  (.I0(\useone/H7[0] ), .I1(\useone/h[0] ), 
            .CI(1'b0), .O(n38), .CO(n39)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i1 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i32  (.I0(\useone/H7[31] ), .I1(\useone/h[31] ), 
            .CI(n863), .O(n861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i31  (.I0(\useone/H7[30] ), .I1(\useone/h[30] ), 
            .CI(n865), .O(n862), .CO(n863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i31 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i30  (.I0(\useone/H7[29] ), .I1(\useone/h[29] ), 
            .CI(n867), .O(n864), .CO(n865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i29  (.I0(\useone/H7[28] ), .I1(\useone/h[28] ), 
            .CI(n869), .O(n866), .CO(n867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i29 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i28  (.I0(\useone/H7[27] ), .I1(\useone/h[27] ), 
            .CI(n871), .O(n868), .CO(n869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i28 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i27  (.I0(\useone/H7[26] ), .I1(\useone/h[26] ), 
            .CI(n873), .O(n870), .CO(n871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i26  (.I0(\useone/H7[25] ), .I1(\useone/h[25] ), 
            .CI(n875), .O(n872), .CO(n873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i26 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i25  (.I0(\useone/H7[24] ), .I1(\useone/h[24] ), 
            .CI(n877), .O(n874), .CO(n875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i25 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i24  (.I0(\useone/H7[23] ), .I1(\useone/h[23] ), 
            .CI(n879), .O(n876), .CO(n877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i24 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i23  (.I0(\useone/H7[22] ), .I1(\useone/h[22] ), 
            .CI(n881), .O(n878), .CO(n879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i23 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i22  (.I0(\useone/H7[21] ), .I1(\useone/h[21] ), 
            .CI(n883), .O(n880), .CO(n881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i22 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i21  (.I0(\useone/H7[20] ), .I1(\useone/h[20] ), 
            .CI(n885), .O(n882), .CO(n883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i20  (.I0(\useone/H7[19] ), .I1(\useone/h[19] ), 
            .CI(n887), .O(n884), .CO(n885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i19  (.I0(\useone/H7[18] ), .I1(\useone/h[18] ), 
            .CI(n889), .O(n886), .CO(n887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i18  (.I0(\useone/H7[17] ), .I1(\useone/h[17] ), 
            .CI(n891), .O(n888), .CO(n889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i17  (.I0(\useone/H7[16] ), .I1(\useone/h[16] ), 
            .CI(n893), .O(n890), .CO(n891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i16  (.I0(\useone/H7[15] ), .I1(\useone/h[15] ), 
            .CI(n895), .O(n892), .CO(n893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i16 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i15  (.I0(\useone/H7[14] ), .I1(\useone/h[14] ), 
            .CI(n897), .O(n894), .CO(n895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i14  (.I0(\useone/H7[13] ), .I1(\useone/h[13] ), 
            .CI(n899), .O(n896), .CO(n897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i13  (.I0(\useone/H7[12] ), .I1(\useone/h[12] ), 
            .CI(n901), .O(n898), .CO(n899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i12  (.I0(\useone/H7[11] ), .I1(\useone/h[11] ), 
            .CI(n903), .O(n900), .CO(n901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i12 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i11  (.I0(\useone/H7[10] ), .I1(\useone/h[10] ), 
            .CI(n905), .O(n902), .CO(n903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i11 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i10  (.I0(\useone/H7[9] ), .I1(\useone/h[9] ), 
            .CI(n907), .O(n904), .CO(n905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i9  (.I0(\useone/H7[8] ), .I1(\useone/h[8] ), 
            .CI(n909), .O(n906), .CO(n907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i9 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i8  (.I0(\useone/H7[7] ), .I1(\useone/h[7] ), 
            .CI(n911), .O(n908), .CO(n909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i7  (.I0(\useone/H7[6] ), .I1(\useone/h[6] ), 
            .CI(n913), .O(n910), .CO(n911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i6  (.I0(\useone/H7[5] ), .I1(\useone/h[5] ), 
            .CI(n915), .O(n912), .CO(n913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i5  (.I0(\useone/H7[4] ), .I1(\useone/h[4] ), 
            .CI(n917), .O(n914), .CO(n915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i5 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i4  (.I0(\useone/H7[3] ), .I1(\useone/h[3] ), 
            .CI(n919), .O(n916), .CO(n917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i4 .I0_POLARITY = 1'b0;
    defparam \useone/add_1022/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1022/i3  (.I0(\useone/H7[2] ), .I1(\useone/h[2] ), 
            .CI(n921), .O(n918), .CO(n919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1022/i2  (.I0(\useone/H7[1] ), .I1(\useone/h[1] ), 
            .CI(n39), .O(n920), .CO(n921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(183)
    defparam \useone/add_1022/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_1022/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i32  (.I0(\useone/H6[31] ), .I1(\useone/g[31] ), 
            .CI(n924), .O(n922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i31  (.I0(\useone/H6[30] ), .I1(\useone/g[30] ), 
            .CI(n926), .O(n923), .CO(n924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i30  (.I0(\useone/H6[29] ), .I1(\useone/g[29] ), 
            .CI(n928), .O(n925), .CO(n926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i29  (.I0(\useone/H6[28] ), .I1(\useone/g[28] ), 
            .CI(n930), .O(n927), .CO(n928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i29 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i28  (.I0(\useone/H6[27] ), .I1(\useone/g[27] ), 
            .CI(n932), .O(n929), .CO(n930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i28 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i27  (.I0(\useone/H6[26] ), .I1(\useone/g[26] ), 
            .CI(n934), .O(n931), .CO(n932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i27 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i26  (.I0(\useone/H6[25] ), .I1(\useone/g[25] ), 
            .CI(n936), .O(n933), .CO(n934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i26 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i25  (.I0(\useone/H6[24] ), .I1(\useone/g[24] ), 
            .CI(n938), .O(n935), .CO(n936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i25 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i24  (.I0(\useone/H6[23] ), .I1(\useone/g[23] ), 
            .CI(n940), .O(n937), .CO(n938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i24 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i24 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i23  (.I0(\useone/H6[22] ), .I1(\useone/g[22] ), 
            .CI(n942), .O(n939), .CO(n940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i22  (.I0(\useone/H6[21] ), .I1(\useone/g[21] ), 
            .CI(n944), .O(n941), .CO(n942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i21  (.I0(\useone/H6[20] ), .I1(\useone/g[20] ), 
            .CI(n946), .O(n943), .CO(n944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i20  (.I0(\useone/H6[19] ), .I1(\useone/g[19] ), 
            .CI(n948), .O(n945), .CO(n946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i19  (.I0(\useone/H6[18] ), .I1(\useone/g[18] ), 
            .CI(n950), .O(n947), .CO(n948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i18  (.I0(\useone/H6[17] ), .I1(\useone/g[17] ), 
            .CI(n952), .O(n949), .CO(n950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i18 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i17  (.I0(\useone/H6[16] ), .I1(\useone/g[16] ), 
            .CI(n954), .O(n951), .CO(n952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i17 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i16  (.I0(\useone/H6[15] ), .I1(\useone/g[15] ), 
            .CI(n956), .O(n953), .CO(n954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i16 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i15  (.I0(\useone/H6[14] ), .I1(\useone/g[14] ), 
            .CI(n958), .O(n955), .CO(n956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i14  (.I0(\useone/H6[13] ), .I1(\useone/g[13] ), 
            .CI(n960), .O(n957), .CO(n958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i13  (.I0(\useone/H6[12] ), .I1(\useone/g[12] ), 
            .CI(n962), .O(n959), .CO(n960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i13 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i12  (.I0(\useone/H6[11] ), .I1(\useone/g[11] ), 
            .CI(n964), .O(n961), .CO(n962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i12 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i11  (.I0(\useone/H6[10] ), .I1(\useone/g[10] ), 
            .CI(n966), .O(n963), .CO(n964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i10  (.I0(\useone/H6[9] ), .I1(\useone/g[9] ), 
            .CI(n968), .O(n965), .CO(n966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i9  (.I0(\useone/H6[8] ), .I1(\useone/g[8] ), 
            .CI(n970), .O(n967), .CO(n968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i9 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i8  (.I0(\useone/H6[7] ), .I1(\useone/g[7] ), 
            .CI(n972), .O(n969), .CO(n970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i8 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i7  (.I0(\useone/H6[6] ), .I1(\useone/g[6] ), 
            .CI(n974), .O(n971), .CO(n972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i6  (.I0(\useone/H6[5] ), .I1(\useone/g[5] ), 
            .CI(n976), .O(n973), .CO(n974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i6 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i5  (.I0(\useone/H6[4] ), .I1(\useone/g[4] ), 
            .CI(n978), .O(n975), .CO(n976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i4  (.I0(\useone/H6[3] ), .I1(\useone/g[3] ), 
            .CI(n980), .O(n977), .CO(n978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i4 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1021/i3  (.I0(\useone/H6[2] ), .I1(\useone/g[2] ), 
            .CI(n982), .O(n979), .CO(n980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1021/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1021/i2  (.I0(\useone/H6[1] ), .I1(\useone/g[1] ), 
            .CI(n37), .O(n981), .CO(n982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(182)
    defparam \useone/add_1021/i2 .I0_POLARITY = 1'b0;
    defparam \useone/add_1021/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i32  (.I0(\useone/H5[31] ), .I1(\useone/f[31] ), 
            .CI(n985), .O(n983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i32 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i31  (.I0(\useone/H5[30] ), .I1(\useone/f[30] ), 
            .CI(n987), .O(n984), .CO(n985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i30  (.I0(\useone/H5[29] ), .I1(\useone/f[29] ), 
            .CI(n989), .O(n986), .CO(n987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i29  (.I0(\useone/H5[28] ), .I1(\useone/f[28] ), 
            .CI(n991), .O(n988), .CO(n989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i29 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i28  (.I0(\useone/H5[27] ), .I1(\useone/f[27] ), 
            .CI(n993), .O(n990), .CO(n991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i28 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i27  (.I0(\useone/H5[26] ), .I1(\useone/f[26] ), 
            .CI(n995), .O(n992), .CO(n993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i26  (.I0(\useone/H5[25] ), .I1(\useone/f[25] ), 
            .CI(n997), .O(n994), .CO(n995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i26 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i25  (.I0(\useone/H5[24] ), .I1(\useone/f[24] ), 
            .CI(n999), .O(n996), .CO(n997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i25 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i24  (.I0(\useone/H5[23] ), .I1(\useone/f[23] ), 
            .CI(n1001), .O(n998), .CO(n999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i23  (.I0(\useone/H5[22] ), .I1(\useone/f[22] ), 
            .CI(n1003), .O(n1000), .CO(n1001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i22  (.I0(\useone/H5[21] ), .I1(\useone/f[21] ), 
            .CI(n1005), .O(n1002), .CO(n1003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i21  (.I0(\useone/H5[20] ), .I1(\useone/f[20] ), 
            .CI(n1007), .O(n1004), .CO(n1005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i20  (.I0(\useone/H5[19] ), .I1(\useone/f[19] ), 
            .CI(n1009), .O(n1006), .CO(n1007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i19  (.I0(\useone/H5[18] ), .I1(\useone/f[18] ), 
            .CI(n1011), .O(n1008), .CO(n1009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i19 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i18  (.I0(\useone/H5[17] ), .I1(\useone/f[17] ), 
            .CI(n1013), .O(n1010), .CO(n1011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i17  (.I0(\useone/H5[16] ), .I1(\useone/f[16] ), 
            .CI(n1015), .O(n1012), .CO(n1013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i17 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i16  (.I0(\useone/H5[15] ), .I1(\useone/f[15] ), 
            .CI(n1017), .O(n1014), .CO(n1015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i16 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i15  (.I0(\useone/H5[14] ), .I1(\useone/f[14] ), 
            .CI(n1019), .O(n1016), .CO(n1017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i14  (.I0(\useone/H5[13] ), .I1(\useone/f[13] ), 
            .CI(n1021), .O(n1018), .CO(n1019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i14 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i13  (.I0(\useone/H5[12] ), .I1(\useone/f[12] ), 
            .CI(n1023), .O(n1020), .CO(n1021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i12  (.I0(\useone/H5[11] ), .I1(\useone/f[11] ), 
            .CI(n1025), .O(n1022), .CO(n1023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i12 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i11  (.I0(\useone/H5[10] ), .I1(\useone/f[10] ), 
            .CI(n1027), .O(n1024), .CO(n1025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i10  (.I0(\useone/H5[9] ), .I1(\useone/f[9] ), 
            .CI(n1029), .O(n1026), .CO(n1027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i9  (.I0(\useone/H5[8] ), .I1(\useone/f[8] ), 
            .CI(n1031), .O(n1028), .CO(n1029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i8  (.I0(\useone/H5[7] ), .I1(\useone/f[7] ), 
            .CI(n1033), .O(n1030), .CO(n1031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i8 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i7  (.I0(\useone/H5[6] ), .I1(\useone/f[6] ), 
            .CI(n1035), .O(n1032), .CO(n1033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i6  (.I0(\useone/H5[5] ), .I1(\useone/f[5] ), 
            .CI(n1037), .O(n1034), .CO(n1035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i5  (.I0(\useone/H5[4] ), .I1(\useone/f[4] ), 
            .CI(n1039), .O(n1036), .CO(n1037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1020/i4  (.I0(\useone/H5[3] ), .I1(\useone/f[3] ), 
            .CI(n1041), .O(n1038), .CO(n1039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i4 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i3  (.I0(\useone/H5[2] ), .I1(\useone/f[2] ), 
            .CI(n1043), .O(n1040), .CO(n1041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i3 .I0_POLARITY = 1'b0;
    defparam \useone/add_1020/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1020/i2  (.I0(\useone/H5[1] ), .I1(\useone/f[1] ), 
            .CI(n35), .O(n1042), .CO(n1043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(181)
    defparam \useone/add_1020/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_1020/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i32  (.I0(\useone/H4[31] ), .I1(\useone/e[31] ), 
            .CI(n1046), .O(n1044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i31  (.I0(\useone/H4[30] ), .I1(\useone/e[30] ), 
            .CI(n1048), .O(n1045), .CO(n1046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i31 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i30  (.I0(\useone/H4[29] ), .I1(\useone/e[29] ), 
            .CI(n1050), .O(n1047), .CO(n1048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i29  (.I0(\useone/H4[28] ), .I1(\useone/e[28] ), 
            .CI(n1052), .O(n1049), .CO(n1050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i29 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i28  (.I0(\useone/H4[27] ), .I1(\useone/e[27] ), 
            .CI(n1054), .O(n1051), .CO(n1052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i28 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i27  (.I0(\useone/H4[26] ), .I1(\useone/e[26] ), 
            .CI(n1056), .O(n1053), .CO(n1054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i26  (.I0(\useone/H4[25] ), .I1(\useone/e[25] ), 
            .CI(n1058), .O(n1055), .CO(n1056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i25  (.I0(\useone/H4[24] ), .I1(\useone/e[24] ), 
            .CI(n1060), .O(n1057), .CO(n1058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i25 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i24  (.I0(\useone/H4[23] ), .I1(\useone/e[23] ), 
            .CI(n1062), .O(n1059), .CO(n1060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i23  (.I0(\useone/H4[22] ), .I1(\useone/e[22] ), 
            .CI(n1064), .O(n1061), .CO(n1062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i22  (.I0(\useone/H4[21] ), .I1(\useone/e[21] ), 
            .CI(n1066), .O(n1063), .CO(n1064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i21  (.I0(\useone/H4[20] ), .I1(\useone/e[20] ), 
            .CI(n1068), .O(n1065), .CO(n1066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i20  (.I0(\useone/H4[19] ), .I1(\useone/e[19] ), 
            .CI(n1070), .O(n1067), .CO(n1068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i20 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i19  (.I0(\useone/H4[18] ), .I1(\useone/e[18] ), 
            .CI(n1072), .O(n1069), .CO(n1070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i19 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i18  (.I0(\useone/H4[17] ), .I1(\useone/e[17] ), 
            .CI(n1074), .O(n1071), .CO(n1072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i18 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i17  (.I0(\useone/H4[16] ), .I1(\useone/e[16] ), 
            .CI(n1076), .O(n1073), .CO(n1074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i16  (.I0(\useone/H4[15] ), .I1(\useone/e[15] ), 
            .CI(n1078), .O(n1075), .CO(n1076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i16 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i15  (.I0(\useone/H4[14] ), .I1(\useone/e[14] ), 
            .CI(n1080), .O(n1077), .CO(n1078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i14  (.I0(\useone/H4[13] ), .I1(\useone/e[13] ), 
            .CI(n1082), .O(n1079), .CO(n1080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i13  (.I0(\useone/H4[12] ), .I1(\useone/e[12] ), 
            .CI(n1084), .O(n1081), .CO(n1082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i13 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i12  (.I0(\useone/H4[11] ), .I1(\useone/e[11] ), 
            .CI(n1086), .O(n1083), .CO(n1084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i11  (.I0(\useone/H4[10] ), .I1(\useone/e[10] ), 
            .CI(n1088), .O(n1085), .CO(n1086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i10  (.I0(\useone/H4[9] ), .I1(\useone/e[9] ), 
            .CI(n1090), .O(n1087), .CO(n1088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i10 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i9  (.I0(\useone/H4[8] ), .I1(\useone/e[8] ), 
            .CI(n1092), .O(n1089), .CO(n1090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i8  (.I0(\useone/H4[7] ), .I1(\useone/e[7] ), 
            .CI(n1094), .O(n1091), .CO(n1092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1019/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1019/i7  (.I0(\useone/H4[6] ), .I1(\useone/e[6] ), 
            .CI(n1096), .O(n1093), .CO(n1094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i7 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i6  (.I0(\useone/H4[5] ), .I1(\useone/e[5] ), 
            .CI(n1098), .O(n1095), .CO(n1096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i6 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i5  (.I0(\useone/H4[4] ), .I1(\useone/e[4] ), 
            .CI(n1100), .O(n1097), .CO(n1098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i5 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i4  (.I0(\useone/H4[3] ), .I1(\useone/e[3] ), 
            .CI(n1102), .O(n1099), .CO(n1100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i4 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i3  (.I0(\useone/H4[2] ), .I1(\useone/e[2] ), 
            .CI(n1104), .O(n1101), .CO(n1102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i3 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1019/i2  (.I0(\useone/H4[1] ), .I1(\useone/e[1] ), 
            .CI(n33), .O(n1103), .CO(n1104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(180)
    defparam \useone/add_1019/i2 .I0_POLARITY = 1'b0;
    defparam \useone/add_1019/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i32  (.I0(\useone/H3[31] ), .I1(\useone/d[31] ), 
            .CI(n1107), .O(n1105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i32 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i31  (.I0(\useone/H3[30] ), .I1(\useone/d[30] ), 
            .CI(n1109), .O(n1106), .CO(n1107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i30  (.I0(\useone/H3[29] ), .I1(\useone/d[29] ), 
            .CI(n1111), .O(n1108), .CO(n1109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i30 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i29  (.I0(\useone/H3[28] ), .I1(\useone/d[28] ), 
            .CI(n1113), .O(n1110), .CO(n1111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i29 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i28  (.I0(\useone/H3[27] ), .I1(\useone/d[27] ), 
            .CI(n1115), .O(n1112), .CO(n1113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i28 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i27  (.I0(\useone/H3[26] ), .I1(\useone/d[26] ), 
            .CI(n1117), .O(n1114), .CO(n1115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i27 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i26  (.I0(\useone/H3[25] ), .I1(\useone/d[25] ), 
            .CI(n1119), .O(n1116), .CO(n1117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i25  (.I0(\useone/H3[24] ), .I1(\useone/d[24] ), 
            .CI(n1121), .O(n1118), .CO(n1119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i25 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i24  (.I0(\useone/H3[23] ), .I1(\useone/d[23] ), 
            .CI(n1123), .O(n1120), .CO(n1121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i23  (.I0(\useone/H3[22] ), .I1(\useone/d[22] ), 
            .CI(n1125), .O(n1122), .CO(n1123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i23 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i22  (.I0(\useone/H3[21] ), .I1(\useone/d[21] ), 
            .CI(n1127), .O(n1124), .CO(n1125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i21  (.I0(\useone/H3[20] ), .I1(\useone/d[20] ), 
            .CI(n1129), .O(n1126), .CO(n1127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i20  (.I0(\useone/H3[19] ), .I1(\useone/d[19] ), 
            .CI(n1131), .O(n1128), .CO(n1129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i20 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i19  (.I0(\useone/H3[18] ), .I1(\useone/d[18] ), 
            .CI(n1133), .O(n1130), .CO(n1131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i19 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i18  (.I0(\useone/H3[17] ), .I1(\useone/d[17] ), 
            .CI(n1135), .O(n1132), .CO(n1133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i18 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i17  (.I0(\useone/H3[16] ), .I1(\useone/d[16] ), 
            .CI(n1137), .O(n1134), .CO(n1135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i17 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i16  (.I0(\useone/H3[15] ), .I1(\useone/d[15] ), 
            .CI(n1139), .O(n1136), .CO(n1137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i16 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i15  (.I0(\useone/H3[14] ), .I1(\useone/d[14] ), 
            .CI(n1141), .O(n1138), .CO(n1139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i14  (.I0(\useone/H3[13] ), .I1(\useone/d[13] ), 
            .CI(n1143), .O(n1140), .CO(n1141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i14 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i13  (.I0(\useone/H3[12] ), .I1(\useone/d[12] ), 
            .CI(n1145), .O(n1142), .CO(n1143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i13 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i12  (.I0(\useone/H3[11] ), .I1(\useone/d[11] ), 
            .CI(n1147), .O(n1144), .CO(n1145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i11  (.I0(\useone/H3[10] ), .I1(\useone/d[10] ), 
            .CI(n1149), .O(n1146), .CO(n1147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i11 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i10  (.I0(\useone/H3[9] ), .I1(\useone/d[9] ), 
            .CI(n1151), .O(n1148), .CO(n1149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i9  (.I0(\useone/H3[8] ), .I1(\useone/d[8] ), 
            .CI(n1153), .O(n1150), .CO(n1151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i9 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i8  (.I0(\useone/H3[7] ), .I1(\useone/d[7] ), 
            .CI(n1155), .O(n1152), .CO(n1153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i7  (.I0(\useone/H3[6] ), .I1(\useone/d[6] ), 
            .CI(n1157), .O(n1154), .CO(n1155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i6  (.I0(\useone/H3[5] ), .I1(\useone/d[5] ), 
            .CI(n1159), .O(n1156), .CO(n1157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i6 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i5  (.I0(\useone/H3[4] ), .I1(\useone/d[4] ), 
            .CI(n1161), .O(n1158), .CO(n1159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i5 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i4  (.I0(\useone/H3[3] ), .I1(\useone/d[3] ), 
            .CI(n1163), .O(n1160), .CO(n1161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i4 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1018/i3  (.I0(\useone/H3[2] ), .I1(\useone/d[2] ), 
            .CI(n1165), .O(n1162), .CO(n1163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1018/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1018/i2  (.I0(\useone/H3[1] ), .I1(\useone/d[1] ), 
            .CI(n31), .O(n1164), .CO(n1165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(179)
    defparam \useone/add_1018/i2 .I0_POLARITY = 1'b0;
    defparam \useone/add_1018/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i32  (.I0(\useone/H2[31] ), .I1(\useone/c[31] ), 
            .CI(n1168), .O(n1166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i31  (.I0(\useone/H2[30] ), .I1(\useone/c[30] ), 
            .CI(n1170), .O(n1167), .CO(n1168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i30  (.I0(\useone/H2[29] ), .I1(\useone/c[29] ), 
            .CI(n1172), .O(n1169), .CO(n1170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i30 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i29  (.I0(\useone/H2[28] ), .I1(\useone/c[28] ), 
            .CI(n1174), .O(n1171), .CO(n1172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i29 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i28  (.I0(\useone/H2[27] ), .I1(\useone/c[27] ), 
            .CI(n1176), .O(n1173), .CO(n1174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i28 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i27  (.I0(\useone/H2[26] ), .I1(\useone/c[26] ), 
            .CI(n1178), .O(n1175), .CO(n1176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i27 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i27 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i26  (.I0(\useone/H2[25] ), .I1(\useone/c[25] ), 
            .CI(n1180), .O(n1177), .CO(n1178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i25  (.I0(\useone/H2[24] ), .I1(\useone/c[24] ), 
            .CI(n1182), .O(n1179), .CO(n1180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i25 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i24  (.I0(\useone/H2[23] ), .I1(\useone/c[23] ), 
            .CI(n1184), .O(n1181), .CO(n1182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i23  (.I0(\useone/H2[22] ), .I1(\useone/c[22] ), 
            .CI(n1186), .O(n1183), .CO(n1184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i23 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i22  (.I0(\useone/H2[21] ), .I1(\useone/c[21] ), 
            .CI(n1188), .O(n1185), .CO(n1186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i22 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i21  (.I0(\useone/H2[20] ), .I1(\useone/c[20] ), 
            .CI(n1190), .O(n1187), .CO(n1188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i20  (.I0(\useone/H2[19] ), .I1(\useone/c[19] ), 
            .CI(n1192), .O(n1189), .CO(n1190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i20 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i19  (.I0(\useone/H2[18] ), .I1(\useone/c[18] ), 
            .CI(n1194), .O(n1191), .CO(n1192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i19 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i18  (.I0(\useone/H2[17] ), .I1(\useone/c[17] ), 
            .CI(n1196), .O(n1193), .CO(n1194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i18 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i17  (.I0(\useone/H2[16] ), .I1(\useone/c[16] ), 
            .CI(n1198), .O(n1195), .CO(n1196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i16  (.I0(\useone/H2[15] ), .I1(\useone/c[15] ), 
            .CI(n1200), .O(n1197), .CO(n1198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i16 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i15  (.I0(\useone/H2[14] ), .I1(\useone/c[14] ), 
            .CI(n1202), .O(n1199), .CO(n1200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i14  (.I0(\useone/H2[13] ), .I1(\useone/c[13] ), 
            .CI(n1204), .O(n1201), .CO(n1202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i14 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i13  (.I0(\useone/H2[12] ), .I1(\useone/c[12] ), 
            .CI(n1206), .O(n1203), .CO(n1204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i13 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i12  (.I0(\useone/H2[11] ), .I1(\useone/c[11] ), 
            .CI(n1208), .O(n1205), .CO(n1206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i11  (.I0(\useone/H2[10] ), .I1(\useone/c[10] ), 
            .CI(n1210), .O(n1207), .CO(n1208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i10  (.I0(\useone/H2[9] ), .I1(\useone/c[9] ), 
            .CI(n1212), .O(n1209), .CO(n1210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i10 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i9  (.I0(\useone/H2[8] ), .I1(\useone/c[8] ), 
            .CI(n1214), .O(n1211), .CO(n1212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i9 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i8  (.I0(\useone/H2[7] ), .I1(\useone/c[7] ), 
            .CI(n1216), .O(n1213), .CO(n1214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i7  (.I0(\useone/H2[6] ), .I1(\useone/c[6] ), 
            .CI(n1218), .O(n1215), .CO(n1216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i7 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i6  (.I0(\useone/H2[5] ), .I1(\useone/c[5] ), 
            .CI(n1220), .O(n1217), .CO(n1218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i6 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i5  (.I0(\useone/H2[4] ), .I1(\useone/c[4] ), 
            .CI(n1222), .O(n1219), .CO(n1220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i5 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1017/i4  (.I0(\useone/H2[3] ), .I1(\useone/c[3] ), 
            .CI(n1224), .O(n1221), .CO(n1222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i4 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i3  (.I0(\useone/H2[2] ), .I1(\useone/c[2] ), 
            .CI(n1226), .O(n1223), .CO(n1224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1017/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1017/i2  (.I0(\useone/H2[1] ), .I1(\useone/c[1] ), 
            .CI(n29), .O(n1225), .CO(n1226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(178)
    defparam \useone/add_1017/i2 .I0_POLARITY = 1'b0;
    defparam \useone/add_1017/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i32  (.I0(\useone/H1[31] ), .I1(\useone/b[31] ), 
            .CI(n1229), .O(n1227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i32 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i32 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i31  (.I0(\useone/H1[30] ), .I1(\useone/b[30] ), 
            .CI(n1231), .O(n1228), .CO(n1229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i30  (.I0(\useone/H1[29] ), .I1(\useone/b[29] ), 
            .CI(n1233), .O(n1230), .CO(n1231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i30 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i29  (.I0(\useone/H1[28] ), .I1(\useone/b[28] ), 
            .CI(n1235), .O(n1232), .CO(n1233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i29 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i29 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i28  (.I0(\useone/H1[27] ), .I1(\useone/b[27] ), 
            .CI(n1237), .O(n1234), .CO(n1235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i28 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i27  (.I0(\useone/H1[26] ), .I1(\useone/b[26] ), 
            .CI(n1239), .O(n1236), .CO(n1237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i26  (.I0(\useone/H1[25] ), .I1(\useone/b[25] ), 
            .CI(n1241), .O(n1238), .CO(n1239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i26 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i25  (.I0(\useone/H1[24] ), .I1(\useone/b[24] ), 
            .CI(n1243), .O(n1240), .CO(n1241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i25 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i25 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i24  (.I0(\useone/H1[23] ), .I1(\useone/b[23] ), 
            .CI(n1245), .O(n1242), .CO(n1243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i23  (.I0(\useone/H1[22] ), .I1(\useone/b[22] ), 
            .CI(n1247), .O(n1244), .CO(n1245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i23 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i23 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i22  (.I0(\useone/H1[21] ), .I1(\useone/b[21] ), 
            .CI(n1249), .O(n1246), .CO(n1247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i22 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i22 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i21  (.I0(\useone/H1[20] ), .I1(\useone/b[20] ), 
            .CI(n1251), .O(n1248), .CO(n1249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i20  (.I0(\useone/H1[19] ), .I1(\useone/b[19] ), 
            .CI(n1253), .O(n1250), .CO(n1251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i19  (.I0(\useone/H1[18] ), .I1(\useone/b[18] ), 
            .CI(n1255), .O(n1252), .CO(n1253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i19 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i19 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i18  (.I0(\useone/H1[17] ), .I1(\useone/b[17] ), 
            .CI(n1257), .O(n1254), .CO(n1255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i18 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i18 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i17  (.I0(\useone/H1[16] ), .I1(\useone/b[16] ), 
            .CI(n1259), .O(n1256), .CO(n1257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i17 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i16  (.I0(\useone/H1[15] ), .I1(\useone/b[15] ), 
            .CI(n1261), .O(n1258), .CO(n1259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i16 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i15  (.I0(\useone/H1[14] ), .I1(\useone/b[14] ), 
            .CI(n1263), .O(n1260), .CO(n1261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i15 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i14  (.I0(\useone/H1[13] ), .I1(\useone/b[13] ), 
            .CI(n1265), .O(n1262), .CO(n1263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i14 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i13  (.I0(\useone/H1[12] ), .I1(\useone/b[12] ), 
            .CI(n1267), .O(n1264), .CO(n1265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i12  (.I0(\useone/H1[11] ), .I1(\useone/b[11] ), 
            .CI(n1269), .O(n1266), .CO(n1267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i12 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i11  (.I0(\useone/H1[10] ), .I1(\useone/b[10] ), 
            .CI(n1271), .O(n1268), .CO(n1269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i11 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i10  (.I0(\useone/H1[9] ), .I1(\useone/b[9] ), 
            .CI(n1273), .O(n1270), .CO(n1271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i10 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i9  (.I0(\useone/H1[8] ), .I1(\useone/b[8] ), 
            .CI(n1275), .O(n1272), .CO(n1273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i8  (.I0(\useone/H1[7] ), .I1(\useone/b[7] ), 
            .CI(n1277), .O(n1274), .CO(n1275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i8 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i7  (.I0(\useone/H1[6] ), .I1(\useone/b[6] ), 
            .CI(n1279), .O(n1276), .CO(n1277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i6  (.I0(\useone/H1[5] ), .I1(\useone/b[5] ), 
            .CI(n1281), .O(n1278), .CO(n1279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i5  (.I0(\useone/H1[4] ), .I1(\useone/b[4] ), 
            .CI(n1283), .O(n1280), .CO(n1281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i4  (.I0(\useone/H1[3] ), .I1(\useone/b[3] ), 
            .CI(n1285), .O(n1282), .CO(n1283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i4 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1016/i3  (.I0(\useone/H1[2] ), .I1(\useone/b[2] ), 
            .CI(n1287), .O(n1284), .CO(n1285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i3 .I0_POLARITY = 1'b0;
    defparam \useone/add_1016/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1016/i2  (.I0(\useone/H1[1] ), .I1(\useone/b[1] ), 
            .CI(n27), .O(n1286), .CO(n1287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(177)
    defparam \useone/add_1016/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_1016/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i32  (.I0(\useone/H0[31] ), .I1(\useone/a[31] ), 
            .CI(n1290), .O(n1288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i31  (.I0(\useone/H0[30] ), .I1(\useone/a[30] ), 
            .CI(n1292), .O(n1289), .CO(n1290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i31 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i31 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i30  (.I0(\useone/H0[29] ), .I1(\useone/a[29] ), 
            .CI(n1294), .O(n1291), .CO(n1292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i30 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i30 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i29  (.I0(\useone/H0[28] ), .I1(\useone/a[28] ), 
            .CI(n1296), .O(n1293), .CO(n1294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i29 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i28  (.I0(\useone/H0[27] ), .I1(\useone/a[27] ), 
            .CI(n1298), .O(n1295), .CO(n1296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i28 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i28 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i27  (.I0(\useone/H0[26] ), .I1(\useone/a[26] ), 
            .CI(n1300), .O(n1297), .CO(n1298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i26  (.I0(\useone/H0[25] ), .I1(\useone/a[25] ), 
            .CI(n1302), .O(n1299), .CO(n1300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i26 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i26 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i25  (.I0(\useone/H0[24] ), .I1(\useone/a[24] ), 
            .CI(n1304), .O(n1301), .CO(n1302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i25 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i24  (.I0(\useone/H0[23] ), .I1(\useone/a[23] ), 
            .CI(n1306), .O(n1303), .CO(n1304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i23  (.I0(\useone/H0[22] ), .I1(\useone/a[22] ), 
            .CI(n1308), .O(n1305), .CO(n1306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i22  (.I0(\useone/H0[21] ), .I1(\useone/a[21] ), 
            .CI(n1310), .O(n1307), .CO(n1308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i21  (.I0(\useone/H0[20] ), .I1(\useone/a[20] ), 
            .CI(n1312), .O(n1309), .CO(n1310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i20  (.I0(\useone/H0[19] ), .I1(\useone/a[19] ), 
            .CI(n1314), .O(n1311), .CO(n1312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i20 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i20 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i19  (.I0(\useone/H0[18] ), .I1(\useone/a[18] ), 
            .CI(n1316), .O(n1313), .CO(n1314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i18  (.I0(\useone/H0[17] ), .I1(\useone/a[17] ), 
            .CI(n1318), .O(n1315), .CO(n1316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i17  (.I0(\useone/H0[16] ), .I1(\useone/a[16] ), 
            .CI(n1320), .O(n1317), .CO(n1318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i17 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i17 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i16  (.I0(\useone/H0[15] ), .I1(\useone/a[15] ), 
            .CI(n1322), .O(n1319), .CO(n1320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i16 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i16 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i15  (.I0(\useone/H0[14] ), .I1(\useone/a[14] ), 
            .CI(n1324), .O(n1321), .CO(n1322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i15 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i14  (.I0(\useone/H0[13] ), .I1(\useone/a[13] ), 
            .CI(n1326), .O(n1323), .CO(n1324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i14 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i14 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i13  (.I0(\useone/H0[12] ), .I1(\useone/a[12] ), 
            .CI(n1328), .O(n1325), .CO(n1326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i12  (.I0(\useone/H0[11] ), .I1(\useone/a[11] ), 
            .CI(n1330), .O(n1327), .CO(n1328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i11  (.I0(\useone/H0[10] ), .I1(\useone/a[10] ), 
            .CI(n1332), .O(n1329), .CO(n1330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i11 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i10  (.I0(\useone/H0[9] ), .I1(\useone/a[9] ), 
            .CI(n1334), .O(n1331), .CO(n1332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i10 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i9  (.I0(\useone/H0[8] ), .I1(\useone/a[8] ), 
            .CI(n1336), .O(n1333), .CO(n1334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i8  (.I0(\useone/H0[7] ), .I1(\useone/a[7] ), 
            .CI(n1338), .O(n1335), .CO(n1336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i7  (.I0(\useone/H0[6] ), .I1(\useone/a[6] ), 
            .CI(n1340), .O(n1337), .CO(n1338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i7 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i6  (.I0(\useone/H0[5] ), .I1(\useone/a[5] ), 
            .CI(n1342), .O(n1339), .CO(n1340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i6 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i5  (.I0(\useone/H0[4] ), .I1(\useone/a[4] ), 
            .CI(n1344), .O(n1341), .CO(n1342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i4  (.I0(\useone/H0[3] ), .I1(\useone/a[3] ), 
            .CI(n1346), .O(n1343), .CO(n1344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i4 .I0_POLARITY = 1'b1;
    defparam \useone/add_1015/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1015/i3  (.I0(\useone/H0[2] ), .I1(\useone/a[2] ), 
            .CI(n1348), .O(n1345), .CO(n1346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i3 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1015/i2  (.I0(\useone/H0[1] ), .I1(\useone/a[1] ), 
            .CI(n25), .O(n1347), .CO(n1348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b0 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(176)
    defparam \useone/add_1015/i2 .I0_POLARITY = 1'b0;
    defparam \useone/add_1015/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \useone/add_1012/i32  (.I0(n1532), .I1(n1471), .CI(n1351), 
            .O(n1349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i31  (.I0(n1533), .I1(n1472), .CI(n1353), 
            .O(n1350), .CO(n1351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i30  (.I0(n1535), .I1(n1474), .CI(n1355), 
            .O(n1352), .CO(n1353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i29  (.I0(n1537), .I1(n1476), .CI(n1357), 
            .O(n1354), .CO(n1355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i29 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i28  (.I0(n1539), .I1(n1478), .CI(n1359), 
            .O(n1356), .CO(n1357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i28 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i27  (.I0(n1541), .I1(n1480), .CI(n1361), 
            .O(n1358), .CO(n1359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i26  (.I0(n1543), .I1(n1482), .CI(n1363), 
            .O(n1360), .CO(n1361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i25  (.I0(n1545), .I1(n1484), .CI(n1365), 
            .O(n1362), .CO(n1363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i25 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i24  (.I0(n1547), .I1(n1486), .CI(n1367), 
            .O(n1364), .CO(n1365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i23  (.I0(n1549), .I1(n1488), .CI(n1369), 
            .O(n1366), .CO(n1367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i22  (.I0(n1551), .I1(n1490), .CI(n1371), 
            .O(n1368), .CO(n1369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i21  (.I0(n1553), .I1(n1492), .CI(n1373), 
            .O(n1370), .CO(n1371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i20  (.I0(n1555), .I1(n1494), .CI(n1375), 
            .O(n1372), .CO(n1373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i19  (.I0(n1557), .I1(n1496), .CI(n1377), 
            .O(n1374), .CO(n1375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i18  (.I0(n1559), .I1(n1498), .CI(n1379), 
            .O(n1376), .CO(n1377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i17  (.I0(n1561), .I1(n1500), .CI(n1381), 
            .O(n1378), .CO(n1379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i16  (.I0(n1563), .I1(n1502), .CI(n1383), 
            .O(n1380), .CO(n1381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i16 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i15  (.I0(n1565), .I1(n1504), .CI(n1385), 
            .O(n1382), .CO(n1383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i15 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i14  (.I0(n1567), .I1(n1506), .CI(n1387), 
            .O(n1384), .CO(n1385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i13  (.I0(n1569), .I1(n1508), .CI(n1389), 
            .O(n1386), .CO(n1387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i12  (.I0(n1571), .I1(n1510), .CI(n1391), 
            .O(n1388), .CO(n1389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i11  (.I0(n1573), .I1(n1512), .CI(n1393), 
            .O(n1390), .CO(n1391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i10  (.I0(n1575), .I1(n1514), .CI(n1395), 
            .O(n1392), .CO(n1393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i9  (.I0(n1577), .I1(n1516), .CI(n1397), 
            .O(n1394), .CO(n1395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i8  (.I0(n1579), .I1(n1518), .CI(n1399), 
            .O(n1396), .CO(n1397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i7  (.I0(n1581), .I1(n1520), .CI(n1401), 
            .O(n1398), .CO(n1399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i6  (.I0(n1583), .I1(n1522), .CI(n1403), 
            .O(n1400), .CO(n1401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i5  (.I0(n1585), .I1(n1524), .CI(n1405), 
            .O(n1402), .CO(n1403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i4  (.I0(n1587), .I1(n1526), .CI(n1407), 
            .O(n1404), .CO(n1405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i4 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i3  (.I0(n1589), .I1(n1528), .CI(n1409), 
            .O(n1406), .CO(n1407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1012/i2  (.I0(n1591), .I1(n1530), .CI(n23), .O(n1408), 
            .CO(n1409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(158)
    defparam \useone/add_1012/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_1012/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i32  (.I0(\useone/d[31] ), .I1(n1532), .CI(n1412), 
            .O(n1410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i32 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i31  (.I0(\useone/d[30] ), .I1(n1533), .CI(n1414), 
            .O(n1411), .CO(n1412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i30  (.I0(\useone/d[29] ), .I1(n1535), .CI(n1416), 
            .O(n1413), .CO(n1414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i30 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i29  (.I0(\useone/d[28] ), .I1(n1537), .CI(n1418), 
            .O(n1415), .CO(n1416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i29 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i28  (.I0(\useone/d[27] ), .I1(n1539), .CI(n1420), 
            .O(n1417), .CO(n1418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i28 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i27  (.I0(\useone/d[26] ), .I1(n1541), .CI(n1422), 
            .O(n1419), .CO(n1420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i27 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i26  (.I0(\useone/d[25] ), .I1(n1543), .CI(n1424), 
            .O(n1421), .CO(n1422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i25  (.I0(\useone/d[24] ), .I1(n1545), .CI(n1426), 
            .O(n1423), .CO(n1424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i25 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i24  (.I0(\useone/d[23] ), .I1(n1547), .CI(n1428), 
            .O(n1425), .CO(n1426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i23  (.I0(\useone/d[22] ), .I1(n1549), .CI(n1430), 
            .O(n1427), .CO(n1428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i23 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i22  (.I0(\useone/d[21] ), .I1(n1551), .CI(n1432), 
            .O(n1429), .CO(n1430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i21  (.I0(\useone/d[20] ), .I1(n1553), .CI(n1434), 
            .O(n1431), .CO(n1432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i20  (.I0(\useone/d[19] ), .I1(n1555), .CI(n1436), 
            .O(n1433), .CO(n1434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i20 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i19  (.I0(\useone/d[18] ), .I1(n1557), .CI(n1438), 
            .O(n1435), .CO(n1436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i19 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i18  (.I0(\useone/d[17] ), .I1(n1559), .CI(n1440), 
            .O(n1437), .CO(n1438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i18 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i17  (.I0(\useone/d[16] ), .I1(n1561), .CI(n1442), 
            .O(n1439), .CO(n1440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i17 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i16  (.I0(\useone/d[15] ), .I1(n1563), .CI(n1444), 
            .O(n1441), .CO(n1442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i16 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i15  (.I0(\useone/d[14] ), .I1(n1565), .CI(n1446), 
            .O(n1443), .CO(n1444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i14  (.I0(\useone/d[13] ), .I1(n1567), .CI(n1448), 
            .O(n1445), .CO(n1446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i14 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i13  (.I0(\useone/d[12] ), .I1(n1569), .CI(n1450), 
            .O(n1447), .CO(n1448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i13 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i12  (.I0(\useone/d[11] ), .I1(n1571), .CI(n1452), 
            .O(n1449), .CO(n1450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i11  (.I0(\useone/d[10] ), .I1(n1573), .CI(n1454), 
            .O(n1451), .CO(n1452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i11 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i10  (.I0(\useone/d[9] ), .I1(n1575), .CI(n1456), 
            .O(n1453), .CO(n1454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i9  (.I0(\useone/d[8] ), .I1(n1577), .CI(n1458), 
            .O(n1455), .CO(n1456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i9 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i8  (.I0(\useone/d[7] ), .I1(n1579), .CI(n1460), 
            .O(n1457), .CO(n1458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i7  (.I0(\useone/d[6] ), .I1(n1581), .CI(n1462), 
            .O(n1459), .CO(n1460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i6  (.I0(\useone/d[5] ), .I1(n1583), .CI(n1464), 
            .O(n1461), .CO(n1462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i6 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i5  (.I0(\useone/d[4] ), .I1(n1585), .CI(n1466), 
            .O(n1463), .CO(n1464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i5 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i4  (.I0(\useone/d[3] ), .I1(n1587), .CI(n1468), 
            .O(n1465), .CO(n1466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i4 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i3  (.I0(\useone/d[2] ), .I1(n1589), .CI(n1470), 
            .O(n1467), .CO(n1468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1011/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1011/i2  (.I0(\useone/d[1] ), .I1(n1591), .CI(n21), 
            .O(n1469), .CO(n1470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(154)
    defparam \useone/add_1011/i2 .I0_POLARITY = 1'b0;
    defparam \useone/add_1011/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i32  (.I0(n3421), .I1(n3422), .CI(n1473), 
            .O(n1471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i31  (.I0(n3424), .I1(n3425), .CI(n1475), 
            .O(n1472), .CO(n1473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i30  (.I0(n3427), .I1(n3428), .CI(n1477), 
            .O(n1474), .CO(n1475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i29  (.I0(n3430), .I1(n3431), .CI(n1479), 
            .O(n1476), .CO(n1477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i29 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i28  (.I0(n3433), .I1(n3434), .CI(n1481), 
            .O(n1478), .CO(n1479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i28 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i27  (.I0(n3436), .I1(n3437), .CI(n1483), 
            .O(n1480), .CO(n1481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i26  (.I0(n3439), .I1(n3440), .CI(n1485), 
            .O(n1482), .CO(n1483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i25  (.I0(n3442), .I1(n3443), .CI(n1487), 
            .O(n1484), .CO(n1485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i25 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i24  (.I0(n3445), .I1(n3446), .CI(n1489), 
            .O(n1486), .CO(n1487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i23  (.I0(n3448), .I1(n3449), .CI(n1491), 
            .O(n1488), .CO(n1489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i22  (.I0(n3451), .I1(n3452), .CI(n1493), 
            .O(n1490), .CO(n1491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i21  (.I0(n3454), .I1(n3455), .CI(n1495), 
            .O(n1492), .CO(n1493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i20  (.I0(n3457), .I1(n3458), .CI(n1497), 
            .O(n1494), .CO(n1495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i19  (.I0(n3460), .I1(n3461), .CI(n1499), 
            .O(n1496), .CO(n1497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i18  (.I0(n3463), .I1(n3464), .CI(n1501), 
            .O(n1498), .CO(n1499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i17  (.I0(n3466), .I1(n3467), .CI(n1503), 
            .O(n1500), .CO(n1501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i16  (.I0(n3469), .I1(n3470), .CI(n1505), 
            .O(n1502), .CO(n1503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i16 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i15  (.I0(n3472), .I1(n3473), .CI(n1507), 
            .O(n1504), .CO(n1505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i15 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i14  (.I0(n3475), .I1(n3476), .CI(n1509), 
            .O(n1506), .CO(n1507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i13  (.I0(n3478), .I1(n3479), .CI(n1511), 
            .O(n1508), .CO(n1509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i12  (.I0(n3481), .I1(n3482), .CI(n1513), 
            .O(n1510), .CO(n1511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i11  (.I0(n3484), .I1(n3485), .CI(n1515), 
            .O(n1512), .CO(n1513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i10  (.I0(n3487), .I1(n3488), .CI(n1517), 
            .O(n1514), .CO(n1515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i9  (.I0(n3490), .I1(n3491), .CI(n1519), 
            .O(n1516), .CO(n1517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i8  (.I0(n3493), .I1(n3494), .CI(n1521), 
            .O(n1518), .CO(n1519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i7  (.I0(n3496), .I1(n3497), .CI(n1523), 
            .O(n1520), .CO(n1521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i6  (.I0(n3499), .I1(n3500), .CI(n1525), 
            .O(n1522), .CO(n1523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i5  (.I0(n3502), .I1(n3503), .CI(n1527), 
            .O(n1524), .CO(n1525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i4  (.I0(n3505), .I1(n3506), .CI(n1529), 
            .O(n1526), .CO(n1527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i4 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i3  (.I0(n3508), .I1(n3509), .CI(n1531), 
            .O(n1528), .CO(n1529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1010/i2  (.I0(n3511), .I1(n3512), .CI(n19), .O(n1530), 
            .CO(n1531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(147)
    defparam \useone/add_1010/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_1010/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i32  (.I0(n1593), .I1(n3515), .CI(n1534), 
            .O(n1532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i31  (.I0(n1594), .I1(n3518), .CI(n1536), 
            .O(n1533), .CO(n1534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i30  (.I0(n1596), .I1(n3521), .CI(n1538), 
            .O(n1535), .CO(n1536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i29  (.I0(n1598), .I1(n3524), .CI(n1540), 
            .O(n1537), .CO(n1538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i29 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i28  (.I0(n1600), .I1(n3527), .CI(n1542), 
            .O(n1539), .CO(n1540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i28 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i27  (.I0(n1602), .I1(n3530), .CI(n1544), 
            .O(n1541), .CO(n1542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i26  (.I0(n1604), .I1(n3533), .CI(n1546), 
            .O(n1543), .CO(n1544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i25  (.I0(n1606), .I1(n3536), .CI(n1548), 
            .O(n1545), .CO(n1546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i25 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i24  (.I0(n1608), .I1(n3539), .CI(n1550), 
            .O(n1547), .CO(n1548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i23  (.I0(n1610), .I1(n3542), .CI(n1552), 
            .O(n1549), .CO(n1550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i22  (.I0(n1612), .I1(n3545), .CI(n1554), 
            .O(n1551), .CO(n1552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i21  (.I0(n1614), .I1(n3548), .CI(n1556), 
            .O(n1553), .CO(n1554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i20  (.I0(n1616), .I1(n3551), .CI(n1558), 
            .O(n1555), .CO(n1556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i19  (.I0(n1618), .I1(n3554), .CI(n1560), 
            .O(n1557), .CO(n1558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i18  (.I0(n1620), .I1(n3557), .CI(n1562), 
            .O(n1559), .CO(n1560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i17  (.I0(n1622), .I1(n3560), .CI(n1564), 
            .O(n1561), .CO(n1562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i16  (.I0(n1624), .I1(n3563), .CI(n1566), 
            .O(n1563), .CO(n1564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i16 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i15  (.I0(n1626), .I1(n3566), .CI(n1568), 
            .O(n1565), .CO(n1566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i15 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i14  (.I0(n1628), .I1(n3569), .CI(n1570), 
            .O(n1567), .CO(n1568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i13  (.I0(n1630), .I1(n3572), .CI(n1572), 
            .O(n1569), .CO(n1570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i12  (.I0(n1632), .I1(n3575), .CI(n1574), 
            .O(n1571), .CO(n1572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i11  (.I0(n1634), .I1(n3578), .CI(n1576), 
            .O(n1573), .CO(n1574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i10  (.I0(n1636), .I1(n3581), .CI(n1578), 
            .O(n1575), .CO(n1576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i9  (.I0(n1638), .I1(n3584), .CI(n1580), 
            .O(n1577), .CO(n1578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i8  (.I0(n1640), .I1(n3587), .CI(n1582), 
            .O(n1579), .CO(n1580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i7  (.I0(n1642), .I1(n3590), .CI(n1584), 
            .O(n1581), .CO(n1582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i6  (.I0(n1644), .I1(n3593), .CI(n1586), 
            .O(n1583), .CO(n1584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i5  (.I0(n1646), .I1(n3596), .CI(n1588), 
            .O(n1585), .CO(n1586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i4  (.I0(n1648), .I1(n3599), .CI(n1590), 
            .O(n1587), .CO(n1588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i4 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i3  (.I0(n1650), .I1(n3602), .CI(n1592), 
            .O(n1589), .CO(n1590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1002/i2  (.I0(n1652), .I1(n3605), .CI(n17), .O(n1591), 
            .CO(n1592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1002/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_1002/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i32  (.I0(n1654), .I1(n3608), .CI(n1595), 
            .O(n1593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i31  (.I0(n1655), .I1(n3611), .CI(n1597), 
            .O(n1594), .CO(n1595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i30  (.I0(n1657), .I1(n3614), .CI(n1599), 
            .O(n1596), .CO(n1597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i29  (.I0(n1659), .I1(n3617), .CI(n1601), 
            .O(n1598), .CO(n1599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i29 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i28  (.I0(n1661), .I1(n3620), .CI(n1603), 
            .O(n1600), .CO(n1601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i28 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i27  (.I0(n1663), .I1(n3623), .CI(n1605), 
            .O(n1602), .CO(n1603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i26  (.I0(n1665), .I1(n3626), .CI(n1607), 
            .O(n1604), .CO(n1605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i25  (.I0(n1667), .I1(n3629), .CI(n1609), 
            .O(n1606), .CO(n1607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i25 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i24  (.I0(n1669), .I1(n3632), .CI(n1611), 
            .O(n1608), .CO(n1609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i23  (.I0(n1671), .I1(n3635), .CI(n1613), 
            .O(n1610), .CO(n1611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i22  (.I0(n1673), .I1(n3638), .CI(n1615), 
            .O(n1612), .CO(n1613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i21  (.I0(n1675), .I1(n3641), .CI(n1617), 
            .O(n1614), .CO(n1615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i20  (.I0(n1677), .I1(n3644), .CI(n1619), 
            .O(n1616), .CO(n1617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i19  (.I0(n1679), .I1(n3647), .CI(n1621), 
            .O(n1618), .CO(n1619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i18  (.I0(n1681), .I1(n3650), .CI(n1623), 
            .O(n1620), .CO(n1621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i17  (.I0(n1683), .I1(n3653), .CI(n1625), 
            .O(n1622), .CO(n1623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i16  (.I0(n1685), .I1(n3656), .CI(n1627), 
            .O(n1624), .CO(n1625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i16 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i15  (.I0(n1687), .I1(n3659), .CI(n1629), 
            .O(n1626), .CO(n1627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i15 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i14  (.I0(n1689), .I1(n3662), .CI(n1631), 
            .O(n1628), .CO(n1629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i13  (.I0(n1691), .I1(n3665), .CI(n1633), 
            .O(n1630), .CO(n1631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i12  (.I0(n1693), .I1(n3668), .CI(n1635), 
            .O(n1632), .CO(n1633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i11  (.I0(n1695), .I1(n3671), .CI(n1637), 
            .O(n1634), .CO(n1635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i10  (.I0(n1697), .I1(n3674), .CI(n1639), 
            .O(n1636), .CO(n1637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i9  (.I0(n1699), .I1(n3677), .CI(n1641), 
            .O(n1638), .CO(n1639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i8  (.I0(n1701), .I1(n3680), .CI(n1643), 
            .O(n1640), .CO(n1641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i7  (.I0(n1703), .I1(n3683), .CI(n1645), 
            .O(n1642), .CO(n1643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i6  (.I0(n1705), .I1(n3686), .CI(n1647), 
            .O(n1644), .CO(n1645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i5  (.I0(n1707), .I1(n3689), .CI(n1649), 
            .O(n1646), .CO(n1647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i4  (.I0(n1709), .I1(n3692), .CI(n1651), 
            .O(n1648), .CO(n1649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i4 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i3  (.I0(n1711), .I1(n3695), .CI(n1653), 
            .O(n1650), .CO(n1651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_1000/i2  (.I0(n1713), .I1(n3698), .CI(n15), .O(n1652), 
            .CO(n1653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_1000/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_1000/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i32  (.I0(n1715), .I1(n3701), .CI(n1656), 
            .O(n1654)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i31  (.I0(n1716), .I1(n3704), .CI(n1658), 
            .O(n1655), .CO(n1656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i31 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i30  (.I0(n1718), .I1(n3707), .CI(n1660), 
            .O(n1657), .CO(n1658)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i29  (.I0(n1720), .I1(n3710), .CI(n1662), 
            .O(n1659), .CO(n1660)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i29 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i28  (.I0(n1722), .I1(n3713), .CI(n1664), 
            .O(n1661), .CO(n1662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i28 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i27  (.I0(n1724), .I1(n3716), .CI(n1666), 
            .O(n1663), .CO(n1664)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i26  (.I0(n1726), .I1(n3719), .CI(n1668), 
            .O(n1665), .CO(n1666)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i26 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i25  (.I0(n1728), .I1(n3722), .CI(n1670), 
            .O(n1667), .CO(n1668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i25 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i24  (.I0(n1730), .I1(n3725), .CI(n1672), 
            .O(n1669), .CO(n1670)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i24 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i23  (.I0(n1732), .I1(n3728), .CI(n1674), 
            .O(n1671), .CO(n1672)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i23 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i22  (.I0(n1734), .I1(n3731), .CI(n1676), 
            .O(n1673), .CO(n1674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i22 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i21  (.I0(n1736), .I1(n3734), .CI(n1678), 
            .O(n1675), .CO(n1676)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i20  (.I0(n1738), .I1(n3737), .CI(n1680), 
            .O(n1677), .CO(n1678)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i19  (.I0(n1740), .I1(n3740), .CI(n1682), 
            .O(n1679), .CO(n1680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i18  (.I0(n1742), .I1(n3743), .CI(n1684), 
            .O(n1681), .CO(n1682)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i17  (.I0(n1744), .I1(n3746), .CI(n1686), 
            .O(n1683), .CO(n1684)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i16  (.I0(n1746), .I1(n3749), .CI(n1688), 
            .O(n1685), .CO(n1686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i16 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i15  (.I0(n1748), .I1(n3752), .CI(n1690), 
            .O(n1687), .CO(n1688)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i15 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i14  (.I0(n1750), .I1(n3755), .CI(n1692), 
            .O(n1689), .CO(n1690)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i13  (.I0(n1752), .I1(n3758), .CI(n1694), 
            .O(n1691), .CO(n1692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i12  (.I0(n1754), .I1(n3761), .CI(n1696), 
            .O(n1693), .CO(n1694)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i12 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i11  (.I0(n1756), .I1(n3764), .CI(n1698), 
            .O(n1695), .CO(n1696)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i11 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i10  (.I0(n1758), .I1(n3767), .CI(n1700), 
            .O(n1697), .CO(n1698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i9  (.I0(n1760), .I1(n3770), .CI(n1702), .O(n1699), 
            .CO(n1700)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i9 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i8  (.I0(n1762), .I1(n3773), .CI(n1704), .O(n1701), 
            .CO(n1702)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i7  (.I0(n1764), .I1(n3776), .CI(n1706), .O(n1703), 
            .CO(n1704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i6  (.I0(n1766), .I1(n3779), .CI(n1708), .O(n1705), 
            .CO(n1706)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i5  (.I0(n1768), .I1(n3782), .CI(n1710), .O(n1707), 
            .CO(n1708)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i5 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i4  (.I0(n1770), .I1(n3785), .CI(n1712), .O(n1709), 
            .CO(n1710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i4 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i3  (.I0(n1772), .I1(n3788), .CI(n1714), .O(n1711), 
            .CO(n1712)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_996/i2  (.I0(n1774), .I1(n3791), .CI(n13), .O(n1713), 
            .CO(n1714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_996/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_996/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i32  (.I0(\useone/h[31] ), .I1(n3793), .CI(n1717), 
            .O(n1715)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i32 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i32 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i31  (.I0(\useone/h[30] ), .I1(n3795), .CI(n1719), 
            .O(n1716), .CO(n1717)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i31 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i31 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i30  (.I0(\useone/h[29] ), .I1(n3797), .CI(n1721), 
            .O(n1718), .CO(n1719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i30 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i30 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i29  (.I0(\useone/h[28] ), .I1(n3799), .CI(n1723), 
            .O(n1720), .CO(n1721)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i29 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i29 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i28  (.I0(\useone/h[27] ), .I1(n3801), .CI(n1725), 
            .O(n1722), .CO(n1723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i28 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i28 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i27  (.I0(\useone/h[26] ), .I1(n3803), .CI(n1727), 
            .O(n1724), .CO(n1725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i27 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i27 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i26  (.I0(\useone/h[25] ), .I1(n3805), .CI(n1729), 
            .O(n1726), .CO(n1727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i26 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i26 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i25  (.I0(\useone/h[24] ), .I1(n3807), .CI(n1731), 
            .O(n1728), .CO(n1729)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i25 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i25 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i24  (.I0(\useone/h[23] ), .I1(n3809), .CI(n1733), 
            .O(n1730), .CO(n1731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i24 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i24 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i23  (.I0(\useone/h[22] ), .I1(n3811), .CI(n1735), 
            .O(n1732), .CO(n1733)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i23 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i23 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i22  (.I0(\useone/h[21] ), .I1(n3813), .CI(n1737), 
            .O(n1734), .CO(n1735)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i22 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i22 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i21  (.I0(\useone/h[20] ), .I1(n3815), .CI(n1739), 
            .O(n1736), .CO(n1737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i21 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i21 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i20  (.I0(\useone/h[19] ), .I1(n3817), .CI(n1741), 
            .O(n1738), .CO(n1739)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i20 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i19  (.I0(\useone/h[18] ), .I1(n3819), .CI(n1743), 
            .O(n1740), .CO(n1741)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i19 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i18  (.I0(\useone/h[17] ), .I1(n3821), .CI(n1745), 
            .O(n1742), .CO(n1743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i18 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i17  (.I0(\useone/h[16] ), .I1(n3823), .CI(n1747), 
            .O(n1744), .CO(n1745)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i17 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i16  (.I0(\useone/h[15] ), .I1(n3825), .CI(n1749), 
            .O(n1746), .CO(n1747)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i16 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i15  (.I0(\useone/h[14] ), .I1(n3827), .CI(n1751), 
            .O(n1748), .CO(n1749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i15 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i14  (.I0(\useone/h[13] ), .I1(n3829), .CI(n1753), 
            .O(n1750), .CO(n1751)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i14 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i13  (.I0(\useone/h[12] ), .I1(n3831), .CI(n1755), 
            .O(n1752), .CO(n1753)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i13 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i12  (.I0(\useone/h[11] ), .I1(n3833), .CI(n1757), 
            .O(n1754), .CO(n1755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i12 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i11  (.I0(\useone/h[10] ), .I1(n3835), .CI(n1759), 
            .O(n1756), .CO(n1757)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i11 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i10  (.I0(\useone/h[9] ), .I1(n3837), .CI(n1761), 
            .O(n1758), .CO(n1759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i10 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i9  (.I0(\useone/h[8] ), .I1(n3839), .CI(n1763), 
            .O(n1760), .CO(n1761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i9 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i8  (.I0(\useone/h[7] ), .I1(n3841), .CI(n1765), 
            .O(n1762), .CO(n1763)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i8 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i7  (.I0(\useone/h[6] ), .I1(n3843), .CI(n1767), 
            .O(n1764), .CO(n1765)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i7 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i6  (.I0(\useone/h[5] ), .I1(n3845), .CI(n1769), 
            .O(n1766), .CO(n1767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i6 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i5  (.I0(\useone/h[4] ), .I1(n3847), .CI(n1771), 
            .O(n1768), .CO(n1769)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i5 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i4  (.I0(\useone/h[3] ), .I1(n3849), .CI(n1773), 
            .O(n1770), .CO(n1771)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b0, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i4 .I0_POLARITY = 1'b0;
    defparam \useone/add_995/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i3  (.I0(\useone/h[2] ), .I1(n3851), .CI(n1775), 
            .O(n1772), .CO(n1773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i3 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \useone/add_995/i2  (.I0(\useone/h[1] ), .I1(n3853), .CI(n11), 
            .O(n1774), .CO(n1775)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // E:\vicharak\effinity_projects\sha_uart\sha_256_fsm_v1.sv(144)
    defparam \useone/add_995/i2 .I0_POLARITY = 1'b1;
    defparam \useone/add_995/i2 .I1_POLARITY = 1'b1;
    EFX_LUT4 LUT__5633 (.I0(\state[0] ), .I1(o_Tx_active), .I2(\state[1] ), 
            .O(ceg_net86)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdbd */ ;
    defparam LUT__5633.LUTMASK = 16'hbdbd;
    EFX_LUT4 LUT__5634 (.I0(\state[0] ), .I1(rst), .I2(hashdone), .I3(\state[1] ), 
            .O(n869_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__5634.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__5635 (.I0(rst), .I1(\state[0] ), .I2(hashdone), .O(n3857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__5635.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__5636 (.I0(\state[0] ), .I1(n3857), .I2(o_Tx_active), 
            .I3(\state[1] ), .O(ceg_net99)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hafec */ ;
    defparam LUT__5636.LUTMASK = 16'hafec;
    EFX_LUT4 LUT__5637 (.I0(\chunk_index[4] ), .I1(\chunk_index[3] ), .I2(\chunk_index[2] ), 
            .O(n3858)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5637.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5638 (.I0(\signature[112] ), .I1(\signature[96] ), .I2(\chunk_index[1] ), 
            .I3(n3858), .O(n3859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__5638.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__5639 (.I0(\chunk_index[3] ), .I1(\chunk_index[2] ), .I2(\chunk_index[4] ), 
            .O(n3860)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5639.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5640 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .I2(\signature[32] ), 
            .I3(\chunk_index[2] ), .O(n3861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5640.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5641 (.I0(n3860), .I1(\signature[160] ), .I2(n3861), 
            .I3(\chunk_index[1] ), .O(n3862)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__5641.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__5642 (.I0(\signature[184] ), .I1(\signature[168] ), .I2(\chunk_index[1] ), 
            .O(n3863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5642.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5643 (.I0(\signature[104] ), .I1(\signature[72] ), .I2(\chunk_index[2] ), 
            .O(n3864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__5643.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__5644 (.I0(\chunk_index[1] ), .I1(\chunk_index[4] ), .I2(\chunk_index[3] ), 
            .O(n3865)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5644.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5645 (.I0(n3864), .I1(n3865), .I2(n3863), .I3(n3860), 
            .O(n3866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__5645.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__5646 (.I0(n3862), .I1(n3859), .I2(n3866), .I3(\chunk_index[0] ), 
            .O(n3867)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fee */ ;
    defparam LUT__5646.LUTMASK = 16'h0fee;
    EFX_LUT4 LUT__5647 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .O(n3868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5647.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5648 (.I0(\signature[216] ), .I1(\signature[200] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n3869)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__5648.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__5649 (.I0(\chunk_index[2] ), .I1(\chunk_index[3] ), .I2(\chunk_index[4] ), 
            .O(n3870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5649.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5650 (.I0(n3868), .I1(\signature[192] ), .I2(n3869), 
            .I3(n3870), .O(n3871)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__5650.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__5651 (.I0(\chunk_index[2] ), .I1(\chunk_index[3] ), .I2(\chunk_index[4] ), 
            .O(n3872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5651.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5652 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .I2(\signature[40] ), 
            .I3(\chunk_index[2] ), .O(n3873)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5652.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5653 (.I0(\chunk_index[1] ), .I1(\chunk_index[0] ), .O(n3874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5653.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5654 (.I0(n3872), .I1(\signature[136] ), .I2(n3873), 
            .I3(n3874), .O(n3875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__5654.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__5655 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .I2(\signature[48] ), 
            .I3(\chunk_index[2] ), .O(n3876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5655.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5656 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .O(n3877)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5656.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5657 (.I0(n3860), .I1(\signature[176] ), .I2(n3876), 
            .I3(n3877), .O(n3878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__5657.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__5658 (.I0(\chunk_index[4] ), .I1(\chunk_index[2] ), .I2(\signature[56] ), 
            .O(n3879)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5658.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5659 (.I0(\signature[152] ), .I1(\signature[24] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[4] ), .O(n3880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__5659.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__5660 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .O(n3881)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5660.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5661 (.I0(n3880), .I1(n3879), .I2(\chunk_index[3] ), 
            .I3(n3881), .O(n3882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__5661.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__5662 (.I0(n3871), .I1(n3875), .I2(n3878), .I3(n3882), 
            .O(n3883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__5662.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__5663 (.I0(\signature[144] ), .I1(\signature[16] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n3884)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__5663.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__5664 (.I0(\signature[240] ), .I1(\signature[80] ), .I2(\chunk_index[2] ), 
            .O(n3885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__5664.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__5665 (.I0(n3885), .I1(n3884), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[3] ), .O(n3886)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hebfc */ ;
    defparam LUT__5665.LUTMASK = 16'hebfc;
    EFX_LUT4 LUT__5666 (.I0(\chunk_index[2] ), .I1(\chunk_index[4] ), .I2(\chunk_index[3] ), 
            .I3(\signature[88] ), .O(n3887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5666.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5667 (.I0(n3858), .I1(\signature[120] ), .I2(n3887), 
            .I3(n3881), .O(n3888)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__5667.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__5668 (.I0(\chunk_index[2] ), .I1(\chunk_index[3] ), .I2(\chunk_index[4] ), 
            .O(n3889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__5668.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__5669 (.I0(\signature[0] ), .I1(\signature[8] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n3890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__5669.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__5670 (.I0(\signature[224] ), .I1(\signature[64] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[4] ), .O(n3891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ff3 */ ;
    defparam LUT__5670.LUTMASK = 16'h5ff3;
    EFX_LUT4 LUT__5671 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\chunk_index[3] ), 
            .O(n3892)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5671.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5672 (.I0(n3891), .I1(n3892), .I2(n3889), .I3(n3890), 
            .O(n3893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__5672.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__5673 (.I0(n3877), .I1(n3886), .I2(n3888), .I3(n3893), 
            .O(n3894)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__5673.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__5674 (.I0(n3872), .I1(n3868), .O(n3895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5674.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5675 (.I0(n3877), .I1(n3870), .I2(\signature[208] ), 
            .O(n3896)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__5675.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__5676 (.I0(\chunk_index[0] ), .I1(\chunk_index[2] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n3897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__5676.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__5677 (.I0(\signature[248] ), .I1(\signature[232] ), .I2(\chunk_index[1] ), 
            .I3(n3897), .O(n3898)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__5677.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__5678 (.I0(\signature[128] ), .I1(n3895), .I2(n3896), 
            .I3(n3898), .O(n3899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__5678.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__5679 (.I0(n3867), .I1(n3883), .I2(n3894), .I3(n3899), 
            .O(n828_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__5679.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__5680 (.I0(\useone/e[6] ), .I1(\useone/e[11] ), .I2(\useone/e[25] ), 
            .O(n1790)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__5680.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__5681 (.I0(\useone/f[0] ), .I1(\useone/g[0] ), .I2(\useone/e[0] ), 
            .O(n1792)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__5681.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__5682 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .O(n3900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5682.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5683 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[6] ), .I3(\useone/round_flag[3] ), .O(n3901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__5683.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__5684 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[2] ), 
            .O(n3902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5684.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5685 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[5] ), .I3(\useone/round_flag[4] ), .O(n3903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5685.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5686 (.I0(n3902), .I1(n3903), .O(n3904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5686.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5687 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[5] ), .O(n3905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5687.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5688 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[3] ), .O(n3906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__5688.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__5689 (.I0(n3905), .I1(n3906), .O(n3907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5689.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5690 (.I0(n3901), .I1(n3900), .I2(n3904), .I3(n3907), 
            .O(n3908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__5690.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__5691 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .O(n3909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5691.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5692 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[3] ), 
            .O(n3910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5692.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5693 (.I0(n3909), .I1(n3910), .O(n3911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5693.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5694 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[6] ), .O(n3912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__5694.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__5695 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .O(n3913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5695.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5696 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[0] ), .O(n3914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5696.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5697 (.I0(n3913), .I1(n3901), .I2(n3903), .I3(n3914), 
            .O(n3915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f */ ;
    defparam LUT__5697.LUTMASK = 16'h035f;
    EFX_LUT4 LUT__5698 (.I0(n3912), .I1(n3911), .I2(n3915), .O(n3916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__5698.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__5699 (.I0(\useone/round_flag[6] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[5] ), .I3(\useone/round_flag[3] ), .O(n3917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__5699.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__5700 (.I0(\useone/round_flag[5] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[4] ), .O(n3918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5700.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5701 (.I0(n3909), .I1(n3917), .I2(n3918), .I3(\useone/round_flag[2] ), 
            .O(n3919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f57 */ ;
    defparam LUT__5701.LUTMASK = 16'h0f57;
    EFX_LUT4 LUT__5702 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[3] ), 
            .O(n3920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5702.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5703 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[0] ), .O(n3921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5703.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5704 (.I0(n3920), .I1(n3921), .O(n3922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5704.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5705 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[5] ), .I3(\useone/round_flag[3] ), .O(n3923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__5705.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__5706 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[6] ), .I3(\useone/round_flag[4] ), .O(n3924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__5706.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__5707 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .O(n3925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5707.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5708 (.I0(n3924), .I1(n3923), .I2(n3925), .O(n3926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__5708.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__5709 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[5] ), .I3(\useone/round_flag[6] ), .O(n3927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__5709.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__5710 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .O(n3928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5710.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5711 (.I0(n3927), .I1(n3917), .I2(n3928), .I3(\useone/round_flag[2] ), 
            .O(n3929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__5711.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__5712 (.I0(n3922), .I1(n3926), .I2(n3929), .I3(n3919), 
            .O(n3930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__5712.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__5713 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .O(n3931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5713.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5714 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .O(n3932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5714.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5715 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[6] ), .I3(\useone/round_flag[5] ), .O(n3933)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__5715.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__5716 (.I0(n3932), .I1(n3931), .I2(n3933), .O(n3934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__5716.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__5717 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .O(n3935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5717.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5718 (.I0(n3917), .I1(n3935), .I2(n3918), .I3(n3914), 
            .O(n3936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__5718.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__5719 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[1] ), 
            .O(n3937)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5719.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5720 (.I0(n3923), .I1(n3900), .I2(n3937), .I3(n3927), 
            .O(n3938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__5720.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__5721 (.I0(n3934), .I1(n3936), .I2(n3938), .O(n3939)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5721.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5722 (.I0(n3908), .I1(n3916), .I2(n3930), .I3(n3939), 
            .O(n1794)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__5722.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__5723 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n3940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f30 */ ;
    defparam LUT__5723.LUTMASK = 16'h1f30;
    EFX_LUT4 LUT__5724 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[1] ), .I3(n3940), .O(n3941)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h55e3 */ ;
    defparam LUT__5724.LUTMASK = 16'h55e3;
    EFX_LUT4 LUT__5725 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[5] ), .O(n3942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb00 */ ;
    defparam LUT__5725.LUTMASK = 16'heb00;
    EFX_LUT4 LUT__5726 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[2] ), 
            .O(n3943)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5726.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5727 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[3] ), 
            .O(n3944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5727.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5728 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .O(n3945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5728.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5729 (.I0(n3943), .I1(n3944), .I2(n3945), .O(n3946)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__5729.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__5730 (.I0(\useone/round_flag[4] ), .I1(n3946), .I2(n3911), 
            .I3(\useone/round_flag[5] ), .O(n3947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__5730.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__5731 (.I0(\useone/state[1] ), .I1(\useone/state[2] ), 
            .I2(\useone/state[0] ), .I3(\i131/useone/w[17][23] ), .O(n1191_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff10 */ ;
    defparam LUT__5731.LUTMASK = 16'hff10;
    EFX_LUT4 LUT__5732 (.I0(n3942), .I1(n3941), .I2(n3947), .I3(n1191_2), 
            .O(n1796)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__5732.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__5733 (.I0(\useone/a[2] ), .I1(\useone/a[13] ), .I2(\useone/a[22] ), 
            .O(n1797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__5733.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__5734 (.I0(\useone/a[0] ), .I1(\useone/b[0] ), .I2(\useone/c[0] ), 
            .O(n1798)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__5734.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__5735 (.I0(rst), .I1(\useone/state[0] ), .I2(\useone/state[1] ), 
            .I3(\useone/state[2] ), .O(\useone/select_1072/Select_0/n5 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__5735.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__5736 (.I0(\useone/state[0] ), .I1(\useone/state[2] ), 
            .I2(\useone/state[1] ), .O(n3948)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__5736.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__5737 (.I0(\useone/round_flag[6] ), .I1(n3948), .I2(\i131/useone/w[17][23] ), 
            .O(\useone/n144202 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__5737.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__5738 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .O(n3949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__5738.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__5739 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[5] ), 
            .O(n3950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5739.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5740 (.I0(\useone/round_flag[4] ), .I1(n3949), .I2(n3950), 
            .I3(\useone/round_flag[6] ), .O(n3951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__5740.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__5741 (.I0(n3951), .I1(n3948), .O(\useone/select_1072/Select_2/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5741.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5742 (.I0(\useone/state[0] ), .I1(\useone/state[1] ), 
            .I2(\useone/state[2] ), .O(\useone/equal_1069/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__5742.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__5743 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[0] ), 
            .O(\useone/select_1071/Select_0/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5743.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5744 (.I0(\useone/state[1] ), .I1(\useone/state[2] ), 
            .I2(\useone/state[0] ), .O(\useone/equal_1067/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__5744.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__5745 (.I0(n3951), .I1(n3948), .I2(\useone/equal_1067/n7 ), 
            .O(\useone/select_1072/Select_1/n8 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__5745.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__5746 (.I0(\useone/select_1072/Select_2/n3 ), .I1(\useone/equal_1069/n7 ), 
            .O(\useone/n39302 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__5746.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__5747 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .O(\useone/n46233 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__5747.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__5748 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .O(n3952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__5748.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__5749 (.I0(n3914), .I1(n3952), .O(\useone/n46238 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__5749.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__5750 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .O(n3953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__5750.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__5751 (.I0(n3953), .I1(\useone/round_flag[3] ), .O(\useone/n46243 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__5751.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__5752 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[3] ), 
            .O(n3954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5752.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5753 (.I0(n3931), .I1(n3954), .O(n3955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5753.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__5754 (.I0(n3955), .I1(\useone/round_flag[4] ), .O(\useone/n46248 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__5754.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__5755 (.I0(n3955), .I1(\useone/round_flag[4] ), .I2(\useone/round_flag[5] ), 
            .O(\useone/n46253 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__5755.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__5756 (.I0(n3955), .I1(\useone/round_flag[4] ), .I2(\useone/round_flag[5] ), 
            .I3(\useone/round_flag[6] ), .O(\useone/n46258 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__5756.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__5757 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[1] ), 
            .O(\useone/select_1071/Select_1/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5757.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5758 (.I0(rst), .I1(\useone/state[0] ), .I2(\useone/state[2] ), 
            .I3(\useone/state[1] ), .O(n3956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h030d */ ;
    defparam LUT__5758.LUTMASK = 16'h030d;
    EFX_LUT4 LUT__5759 (.I0(n3956), .I1(\signature[2] ), .I2(\useone/equal_1069/n7 ), 
            .I3(\useone/H7[2] ), .O(\useone/n39297 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__5759.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__5760 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[3] ), 
            .O(\useone/select_1071/Select_3/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5760.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5761 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[4] ), 
            .O(\useone/select_1071/Select_4/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5761.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5762 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[5] ), 
            .O(\useone/select_1071/Select_5/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5762.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5763 (.I0(n3956), .I1(\signature[6] ), .I2(\useone/equal_1069/n7 ), 
            .I3(\useone/H7[6] ), .O(\useone/n39293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__5763.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__5764 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[7] ), 
            .O(\useone/select_1071/Select_7/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5764.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5765 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[8] ), 
            .O(\useone/select_1071/Select_8/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5765.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5766 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[9] ), 
            .O(\useone/select_1071/Select_9/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5766.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5767 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[10] ), 
            .O(\useone/select_1071/Select_10/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5767.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5768 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[11] ), 
            .O(\useone/select_1071/Select_11/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5768.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5769 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[12] ), 
            .O(\useone/select_1071/Select_12/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5769.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5770 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[13] ), 
            .O(\useone/select_1071/Select_13/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5770.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5771 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[14] ), 
            .O(\useone/select_1071/Select_14/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5771.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5772 (.I0(n3956), .I1(\signature[15] ), .I2(\useone/equal_1069/n7 ), 
            .I3(\useone/H7[15] ), .O(\useone/n39284 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h888f */ ;
    defparam LUT__5772.LUTMASK = 16'h888f;
    EFX_LUT4 LUT__5773 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[16] ), 
            .O(\useone/select_1071/Select_16/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5773.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5774 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[17] ), 
            .O(\useone/select_1071/Select_17/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5774.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5775 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[18] ), 
            .O(\useone/select_1071/Select_18/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5775.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5776 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[19] ), 
            .O(\useone/select_1071/Select_19/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5776.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5777 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[20] ), 
            .O(\useone/select_1071/Select_20/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5777.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5778 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[21] ), 
            .O(\useone/select_1071/Select_21/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5778.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5779 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[22] ), 
            .O(\useone/select_1071/Select_22/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5779.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5780 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[23] ), 
            .O(\useone/select_1071/Select_23/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5780.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5781 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[24] ), 
            .O(\useone/select_1071/Select_24/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5781.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5782 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[25] ), 
            .O(\useone/select_1071/Select_25/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5782.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5783 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[26] ), 
            .O(\useone/select_1071/Select_26/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5783.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5784 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[27] ), 
            .O(\useone/select_1071/Select_27/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5784.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5785 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[28] ), 
            .O(\useone/select_1071/Select_28/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5785.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5786 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[29] ), 
            .O(\useone/select_1071/Select_29/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5786.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5787 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[30] ), 
            .O(\useone/select_1071/Select_30/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5787.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5788 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H7[31] ), 
            .O(\useone/select_1071/Select_31/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5788.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5789 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[0] ), 
            .O(\useone/select_1071/Select_32/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5789.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5790 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[1] ), 
            .O(\useone/select_1071/Select_33/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5790.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5791 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[2] ), 
            .O(\useone/select_1071/Select_34/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5791.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5792 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[3] ), 
            .O(\useone/select_1071/Select_35/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5792.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5793 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[4] ), 
            .O(\useone/select_1071/Select_36/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5793.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5794 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[5] ), 
            .O(\useone/select_1071/Select_37/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5794.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5795 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[6] ), 
            .O(\useone/select_1071/Select_38/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5795.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5796 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[7] ), 
            .O(\useone/select_1071/Select_39/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5796.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5797 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[8] ), 
            .O(\useone/select_1071/Select_40/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5797.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5798 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[9] ), 
            .O(\useone/select_1071/Select_41/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5798.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5799 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[10] ), 
            .O(\useone/select_1071/Select_42/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5799.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5800 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[11] ), 
            .O(\useone/select_1071/Select_43/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5800.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5801 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[12] ), 
            .O(\useone/select_1071/Select_44/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5801.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5802 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[13] ), 
            .O(\useone/select_1071/Select_45/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5802.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5803 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[14] ), 
            .O(\useone/select_1071/Select_46/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5803.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5804 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[15] ), 
            .O(\useone/select_1071/Select_47/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5804.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5805 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[16] ), 
            .O(\useone/select_1071/Select_48/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5805.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5806 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[17] ), 
            .O(\useone/select_1071/Select_49/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5806.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5807 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[18] ), 
            .O(\useone/select_1071/Select_50/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5807.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5808 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[19] ), 
            .O(\useone/select_1071/Select_51/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5808.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5809 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[20] ), 
            .O(\useone/select_1071/Select_52/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5809.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5810 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[21] ), 
            .O(\useone/select_1071/Select_53/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5810.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5811 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[22] ), 
            .O(\useone/select_1071/Select_54/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5811.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5812 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[23] ), 
            .O(\useone/select_1071/Select_55/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5812.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5813 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[24] ), 
            .O(\useone/select_1071/Select_56/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5813.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5814 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[25] ), 
            .O(\useone/select_1071/Select_57/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5814.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5815 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[26] ), 
            .O(\useone/select_1071/Select_58/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5815.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5816 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[27] ), 
            .O(\useone/select_1071/Select_59/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5816.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5817 (.I0(\useone/H6[28] ), .I1(\useone/equal_1069/n7 ), 
            .I2(n3948), .I3(\signature[60] ), .O(\useone/n39239 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf111 */ ;
    defparam LUT__5817.LUTMASK = 16'hf111;
    EFX_LUT4 LUT__5818 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[29] ), 
            .O(\useone/select_1071/Select_61/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5818.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5819 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[30] ), 
            .O(\useone/select_1071/Select_62/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5819.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5820 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H6[31] ), 
            .O(\useone/select_1071/Select_63/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5820.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5821 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[0] ), 
            .O(\useone/select_1071/Select_64/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5821.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5822 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[1] ), 
            .O(\useone/select_1071/Select_65/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5822.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5823 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[2] ), 
            .O(\useone/select_1071/Select_66/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5823.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5824 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[3] ), 
            .O(\useone/select_1071/Select_67/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5824.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5825 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[4] ), 
            .O(\useone/select_1071/Select_68/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5825.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5826 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[5] ), 
            .O(\useone/select_1071/Select_69/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5826.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5827 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[6] ), 
            .O(\useone/select_1071/Select_70/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5827.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5828 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[7] ), 
            .O(\useone/select_1071/Select_71/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5828.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5829 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[8] ), 
            .O(\useone/select_1071/Select_72/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5829.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5830 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[9] ), 
            .O(\useone/select_1071/Select_73/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5830.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5831 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[10] ), 
            .O(\useone/select_1071/Select_74/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5831.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5832 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[11] ), 
            .O(\useone/select_1071/Select_75/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5832.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5833 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[12] ), 
            .O(\useone/select_1071/Select_76/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5833.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5834 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[13] ), 
            .O(\useone/select_1071/Select_77/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5834.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5835 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[14] ), 
            .O(\useone/select_1071/Select_78/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5835.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5836 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[15] ), 
            .O(\useone/select_1071/Select_79/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5836.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5837 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[16] ), 
            .O(\useone/select_1071/Select_80/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5837.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5838 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[17] ), 
            .O(\useone/select_1071/Select_81/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5838.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5839 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[18] ), 
            .O(\useone/select_1071/Select_82/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5839.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5840 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[19] ), 
            .O(\useone/select_1071/Select_83/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5840.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5841 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[20] ), 
            .O(\useone/select_1071/Select_84/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5841.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5842 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[21] ), 
            .O(\useone/select_1071/Select_85/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5842.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5843 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[22] ), 
            .O(\useone/select_1071/Select_86/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5843.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5844 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[23] ), 
            .O(\useone/select_1071/Select_87/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5844.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5845 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[24] ), 
            .O(\useone/select_1071/Select_88/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5845.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5846 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[25] ), 
            .O(\useone/select_1071/Select_89/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5846.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5847 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[26] ), 
            .O(\useone/select_1071/Select_90/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5847.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5848 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[27] ), 
            .O(\useone/select_1071/Select_91/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5848.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5849 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[28] ), 
            .O(\useone/select_1071/Select_92/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5849.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5850 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[29] ), 
            .O(\useone/select_1071/Select_93/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5850.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5851 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[30] ), 
            .O(\useone/select_1071/Select_94/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5851.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5852 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H5[31] ), 
            .O(\useone/select_1071/Select_95/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5852.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5853 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[0] ), 
            .O(\useone/select_1071/Select_96/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5853.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5854 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[1] ), 
            .O(\useone/select_1071/Select_97/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5854.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5855 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[2] ), 
            .O(\useone/select_1071/Select_98/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5855.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5856 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[3] ), 
            .O(\useone/select_1071/Select_99/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5856.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5857 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[4] ), 
            .O(\useone/select_1071/Select_100/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5857.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5858 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[5] ), 
            .O(\useone/select_1071/Select_101/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5858.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5859 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[6] ), 
            .O(\useone/select_1071/Select_102/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5859.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5860 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[7] ), 
            .O(\useone/select_1071/Select_103/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5860.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5861 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[8] ), 
            .O(\useone/select_1071/Select_104/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5861.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5862 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[9] ), 
            .O(\useone/select_1071/Select_105/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5862.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5863 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[10] ), 
            .O(\useone/select_1071/Select_106/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5863.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5864 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[11] ), 
            .O(\useone/select_1071/Select_107/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5864.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5865 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[12] ), 
            .O(\useone/select_1071/Select_108/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5865.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5866 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[13] ), 
            .O(\useone/select_1071/Select_109/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5866.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5867 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[14] ), 
            .O(\useone/select_1071/Select_110/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5867.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5868 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[15] ), 
            .O(\useone/select_1071/Select_111/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5868.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5869 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[16] ), 
            .O(\useone/select_1071/Select_112/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5869.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5870 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[17] ), 
            .O(\useone/select_1071/Select_113/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5870.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5871 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[18] ), 
            .O(\useone/select_1071/Select_114/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5871.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5872 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[19] ), 
            .O(\useone/select_1071/Select_115/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5872.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5873 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[20] ), 
            .O(\useone/select_1071/Select_116/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5873.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5874 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[21] ), 
            .O(\useone/select_1071/Select_117/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5874.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5875 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[22] ), 
            .O(\useone/select_1071/Select_118/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5875.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5876 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[23] ), 
            .O(\useone/select_1071/Select_119/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5876.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5877 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[24] ), 
            .O(\useone/select_1071/Select_120/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5877.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5878 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[25] ), 
            .O(\useone/select_1071/Select_121/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5878.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5879 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[26] ), 
            .O(\useone/select_1071/Select_122/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5879.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5880 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[27] ), 
            .O(\useone/select_1071/Select_123/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5880.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5881 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[28] ), 
            .O(\useone/select_1071/Select_124/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5881.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5882 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[29] ), 
            .O(\useone/select_1071/Select_125/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5882.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5883 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[30] ), 
            .O(\useone/select_1071/Select_126/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5883.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5884 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H4[31] ), 
            .O(\useone/select_1071/Select_127/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5884.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5885 (.I0(n3956), .I1(\signature[128] ), .I2(\useone/equal_1069/n7 ), 
            .I3(\useone/H3[0] ), .O(\useone/n39171 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f88 */ ;
    defparam LUT__5885.LUTMASK = 16'h8f88;
    EFX_LUT4 LUT__5886 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[1] ), 
            .O(\useone/select_1071/Select_129/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5886.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5887 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[2] ), 
            .O(\useone/select_1071/Select_130/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5887.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5888 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[3] ), 
            .O(\useone/select_1071/Select_131/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5888.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5889 (.I0(\useone/H3[4] ), .I1(\useone/equal_1069/n7 ), 
            .I2(n3948), .I3(\signature[132] ), .O(\useone/n39167 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf111 */ ;
    defparam LUT__5889.LUTMASK = 16'hf111;
    EFX_LUT4 LUT__5890 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[5] ), 
            .O(\useone/select_1071/Select_133/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5890.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5891 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[6] ), 
            .O(\useone/select_1071/Select_134/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5891.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5892 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[7] ), 
            .O(\useone/select_1071/Select_135/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5892.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5893 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[8] ), 
            .O(\useone/select_1071/Select_136/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5893.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5894 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[9] ), 
            .O(\useone/select_1071/Select_137/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5894.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5895 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[10] ), 
            .O(\useone/select_1071/Select_138/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5895.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5896 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[11] ), 
            .O(\useone/select_1071/Select_139/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5896.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5897 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[12] ), 
            .O(\useone/select_1071/Select_140/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5897.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5898 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[13] ), 
            .O(\useone/select_1071/Select_141/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5898.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5899 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[14] ), 
            .O(\useone/select_1071/Select_142/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5899.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5900 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[15] ), 
            .O(\useone/select_1071/Select_143/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5900.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5901 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[16] ), 
            .O(\useone/select_1071/Select_144/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5901.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5902 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[17] ), 
            .O(\useone/select_1071/Select_145/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5902.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5903 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[18] ), 
            .O(\useone/select_1071/Select_146/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5903.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5904 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[19] ), 
            .O(\useone/select_1071/Select_147/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5904.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5905 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[20] ), 
            .O(\useone/select_1071/Select_148/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5905.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5906 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[21] ), 
            .O(\useone/select_1071/Select_149/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5906.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5907 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[22] ), 
            .O(\useone/select_1071/Select_150/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5907.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5908 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[23] ), 
            .O(\useone/select_1071/Select_151/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5908.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5909 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[24] ), 
            .O(\useone/select_1071/Select_152/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5909.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5910 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[25] ), 
            .O(\useone/select_1071/Select_153/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5910.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5911 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[26] ), 
            .O(\useone/select_1071/Select_154/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5911.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5912 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[27] ), 
            .O(\useone/select_1071/Select_155/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5912.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5913 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[28] ), 
            .O(\useone/select_1071/Select_156/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5913.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5914 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[29] ), 
            .O(\useone/select_1071/Select_157/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5914.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5915 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[30] ), 
            .O(\useone/select_1071/Select_158/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5915.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5916 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H3[31] ), 
            .O(\useone/select_1071/Select_159/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5916.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5917 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[0] ), 
            .O(\useone/select_1071/Select_160/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5917.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5918 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[1] ), 
            .O(\useone/select_1071/Select_161/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5918.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5919 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[2] ), 
            .O(\useone/select_1071/Select_162/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5919.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5920 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[3] ), 
            .O(\useone/select_1071/Select_163/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5920.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5921 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[4] ), 
            .O(\useone/select_1071/Select_164/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5921.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5922 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[5] ), 
            .O(\useone/select_1071/Select_165/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5922.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5923 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[6] ), 
            .O(\useone/select_1071/Select_166/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5923.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5924 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[7] ), 
            .O(\useone/select_1071/Select_167/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5924.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5925 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[8] ), 
            .O(\useone/select_1071/Select_168/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5925.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5926 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[9] ), 
            .O(\useone/select_1071/Select_169/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5926.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5927 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[10] ), 
            .O(\useone/select_1071/Select_170/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5927.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5928 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[11] ), 
            .O(\useone/select_1071/Select_171/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5928.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5929 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[12] ), 
            .O(\useone/select_1071/Select_172/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5929.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5930 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[13] ), 
            .O(\useone/select_1071/Select_173/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5930.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5931 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[14] ), 
            .O(\useone/select_1071/Select_174/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5931.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5932 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[15] ), 
            .O(\useone/select_1071/Select_175/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5932.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5933 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[16] ), 
            .O(\useone/select_1071/Select_176/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5933.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5934 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[17] ), 
            .O(\useone/select_1071/Select_177/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5934.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5935 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[18] ), 
            .O(\useone/select_1071/Select_178/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5935.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5936 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[19] ), 
            .O(\useone/select_1071/Select_179/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5936.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5937 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[20] ), 
            .O(\useone/select_1071/Select_180/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5937.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5938 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[21] ), 
            .O(\useone/select_1071/Select_181/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5938.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5939 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[22] ), 
            .O(\useone/select_1071/Select_182/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5939.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5940 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[23] ), 
            .O(\useone/select_1071/Select_183/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5940.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5941 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[24] ), 
            .O(\useone/select_1071/Select_184/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5941.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5942 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[25] ), 
            .O(\useone/select_1071/Select_185/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5942.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5943 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[26] ), 
            .O(\useone/select_1071/Select_186/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5943.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5944 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[27] ), 
            .O(\useone/select_1071/Select_187/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5944.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5945 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[28] ), 
            .O(\useone/select_1071/Select_188/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5945.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5946 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[29] ), 
            .O(\useone/select_1071/Select_189/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5946.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5947 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[30] ), 
            .O(\useone/select_1071/Select_190/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5947.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5948 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H2[31] ), 
            .O(\useone/select_1071/Select_191/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5948.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5949 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[0] ), 
            .O(\useone/select_1071/Select_192/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5949.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5950 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[1] ), 
            .O(\useone/select_1071/Select_193/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5950.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5951 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[2] ), 
            .O(\useone/select_1071/Select_194/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5951.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5952 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[3] ), 
            .O(\useone/select_1071/Select_195/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5952.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5953 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[4] ), 
            .O(\useone/select_1071/Select_196/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5953.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5954 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[5] ), 
            .O(\useone/select_1071/Select_197/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5954.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5955 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[6] ), 
            .O(\useone/select_1071/Select_198/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5955.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5956 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[7] ), 
            .O(\useone/select_1071/Select_199/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5956.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5957 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[8] ), 
            .O(\useone/select_1071/Select_200/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5957.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5958 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[9] ), 
            .O(\useone/select_1071/Select_201/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5958.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5959 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[10] ), 
            .O(\useone/select_1071/Select_202/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5959.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5960 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[11] ), 
            .O(\useone/select_1071/Select_203/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5960.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5961 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[12] ), 
            .O(\useone/select_1071/Select_204/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5961.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5962 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[13] ), 
            .O(\useone/select_1071/Select_205/n6 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5962.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5963 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[14] ), 
            .O(\useone/select_1071/Select_206/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5963.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5964 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[15] ), 
            .O(\useone/select_1071/Select_207/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5964.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5965 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[16] ), 
            .O(\useone/select_1071/Select_208/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5965.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5966 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[17] ), 
            .O(\useone/select_1071/Select_209/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5966.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5967 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[18] ), 
            .O(\useone/select_1071/Select_210/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5967.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5968 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[19] ), 
            .O(\useone/select_1071/Select_211/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5968.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5969 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[20] ), 
            .O(\useone/select_1071/Select_212/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5969.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5970 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[21] ), 
            .O(\useone/select_1071/Select_213/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5970.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5971 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[22] ), 
            .O(\useone/select_1071/Select_214/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5971.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5972 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[23] ), 
            .O(\useone/select_1071/Select_215/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5972.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5973 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[24] ), 
            .O(\useone/select_1071/Select_216/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5973.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5974 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[25] ), 
            .O(\useone/select_1071/Select_217/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5974.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5975 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[26] ), 
            .O(\useone/select_1071/Select_218/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5975.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5976 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[27] ), 
            .O(\useone/select_1071/Select_219/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5976.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5977 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[28] ), 
            .O(\useone/select_1071/Select_220/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5977.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5978 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[29] ), 
            .O(\useone/select_1071/Select_221/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5978.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5979 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[30] ), 
            .O(\useone/select_1071/Select_222/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5979.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5980 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H1[31] ), 
            .O(\useone/select_1071/Select_223/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5980.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5981 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[0] ), 
            .O(\useone/select_1071/Select_224/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5981.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5982 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[1] ), 
            .O(\useone/select_1071/Select_225/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5982.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5983 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[2] ), 
            .O(\useone/select_1071/Select_226/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5983.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5984 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[3] ), 
            .O(\useone/select_1071/Select_227/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5984.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5985 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[4] ), 
            .O(\useone/select_1071/Select_228/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5985.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5986 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[5] ), 
            .O(\useone/select_1071/Select_229/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5986.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5987 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[6] ), 
            .O(\useone/select_1071/Select_230/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5987.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5988 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[7] ), 
            .O(\useone/select_1071/Select_231/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5988.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5989 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[8] ), 
            .O(\useone/select_1071/Select_232/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5989.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5990 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[9] ), 
            .O(\useone/select_1071/Select_233/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5990.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5991 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[10] ), 
            .O(\useone/select_1071/Select_234/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5991.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5992 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[11] ), 
            .O(\useone/select_1071/Select_235/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5992.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5993 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[12] ), 
            .O(\useone/select_1071/Select_236/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5993.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5994 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[13] ), 
            .O(\useone/select_1071/Select_237/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5994.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5995 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[14] ), 
            .O(\useone/select_1071/Select_238/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5995.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5996 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[15] ), 
            .O(\useone/select_1071/Select_239/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5996.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5997 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[16] ), 
            .O(\useone/select_1071/Select_240/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__5997.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__5998 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[17] ), 
            .O(\useone/select_1071/Select_241/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5998.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__5999 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[18] ), 
            .O(\useone/select_1071/Select_242/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__5999.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6000 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[19] ), 
            .O(\useone/select_1071/Select_243/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6000.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6001 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[20] ), 
            .O(\useone/select_1071/Select_244/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6001.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6002 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[21] ), 
            .O(\useone/select_1071/Select_245/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6002.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6003 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[22] ), 
            .O(\useone/select_1071/Select_246/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6003.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6004 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[23] ), 
            .O(\useone/select_1071/Select_247/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6004.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6005 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[24] ), 
            .O(\useone/select_1071/Select_248/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6005.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6006 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[25] ), 
            .O(\useone/select_1071/Select_249/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6006.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6007 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[26] ), 
            .O(\useone/select_1071/Select_250/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6007.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6008 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[27] ), 
            .O(\useone/select_1071/Select_251/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6008.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6009 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[28] ), 
            .O(\useone/select_1071/Select_252/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6009.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6010 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[29] ), 
            .O(\useone/select_1071/Select_253/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6010.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6011 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[30] ), 
            .O(\useone/select_1071/Select_254/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6011.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6012 (.I0(\useone/equal_1069/n7 ), .I1(\useone/H0[31] ), 
            .O(\useone/select_1071/Select_255/n2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6012.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6013 (.I0(\useuart/r_Clock_Count[4] ), .I1(\useuart/r_Clock_Count[3] ), 
            .I2(\useuart/r_Clock_Count[5] ), .I3(\useuart/r_Clock_Count[6] ), 
            .O(n3957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6013.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6014 (.I0(\useuart/r_Clock_Count[7] ), .I1(\useuart/r_Clock_Count[8] ), 
            .I2(\useuart/r_Clock_Count[9] ), .I3(\useuart/r_Clock_Count[11] ), 
            .O(n3958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6014.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6015 (.I0(\useuart/r_Clock_Count[11] ), .I1(\useuart/r_Clock_Count[10] ), 
            .I2(\useuart/r_Clock_Count[12] ), .O(n3959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6015.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6016 (.I0(n3957), .I1(n3958), .I2(n3959), .O(\useuart/LessThan_9/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__6016.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__6017 (.I0(\useuart/r_SM_Main[1] ), .I1(\useuart/r_SM_Main[0] ), 
            .I2(\useuart/LessThan_9/n26 ), .O(n3960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6017.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6018 (.I0(\useuart/r_Clock_Count[0] ), .I1(n3960), .O(\useuart/n844 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6018.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6019 (.I0(\useuart/r_Tx_Data[2] ), .I1(\useuart/r_Tx_Data[0] ), 
            .I2(\useuart/r_Bit_Index[1] ), .O(n3961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6019.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6020 (.I0(\useuart/r_Tx_Data[1] ), .I1(\useuart/r_Tx_Data[3] ), 
            .I2(\useuart/r_Bit_Index[1] ), .O(n3962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6020.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6021 (.I0(n3962), .I1(n3961), .I2(\useuart/r_Bit_Index[2] ), 
            .I3(\useuart/r_Bit_Index[0] ), .O(n3963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0503 */ ;
    defparam LUT__6021.LUTMASK = 16'h0503;
    EFX_LUT4 LUT__6022 (.I0(\useuart/r_Tx_Data[4] ), .I1(\useuart/r_Tx_Data[6] ), 
            .I2(\useuart/r_Bit_Index[1] ), .O(n3964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6022.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6023 (.I0(\useuart/r_Tx_Data[5] ), .I1(\useuart/r_Tx_Data[7] ), 
            .I2(\useuart/r_Bit_Index[1] ), .O(n3965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6023.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6024 (.I0(n3965), .I1(n3964), .I2(\useuart/r_Bit_Index[0] ), 
            .I3(\useuart/r_Bit_Index[2] ), .O(n3966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6024.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6025 (.I0(n3963), .I1(n3966), .I2(\useuart/r_SM_Main[0] ), 
            .I3(\useuart/r_SM_Main[1] ), .O(\useuart/n634 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe0f */ ;
    defparam LUT__6025.LUTMASK = 16'hfe0f;
    EFX_LUT4 LUT__6026 (.I0(\useuart/r_Bit_Index[0] ), .I1(\useuart/r_SM_Main[1] ), 
            .O(\useuart/n848 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6026.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6027 (.I0(\useuart/r_SM_Main[1] ), .I1(\useuart/LessThan_9/n26 ), 
            .I2(\useuart/r_SM_Main[0] ), .I3(\useuart/r_SM_Main[2] ), .O(ceg_net79)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__6027.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__6028 (.I0(\useuart/r_SM_Main[2] ), .I1(\useuart/r_SM_Main[1] ), 
            .I2(\useuart/r_SM_Main[0] ), .O(\useuart/n942 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6028.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6029 (.I0(\useuart/r_SM_Main[1] ), .I1(tx_valid), .O(n3967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6029.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6030 (.I0(\useuart/r_SM_Main[0] ), .I1(\useuart/r_SM_Main[2] ), 
            .I2(n3967), .O(\useuart/n960 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6030.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6031 (.I0(\useuart/n942 ), .I1(\useuart/LessThan_9/n26 ), 
            .I2(\useuart/n960 ), .O(ceg_net77)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6031.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6032 (.I0(\useuart/r_Bit_Index[0] ), .I1(\useuart/r_Bit_Index[1] ), 
            .I2(\useuart/r_Bit_Index[2] ), .I3(\useuart/r_SM_Main[1] ), 
            .O(n3968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6032.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6033 (.I0(n3968), .I1(n3967), .I2(\useuart/LessThan_9/n26 ), 
            .I3(\useuart/r_SM_Main[0] ), .O(\useuart/n840 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ce */ ;
    defparam LUT__6033.LUTMASK = 16'hf0ce;
    EFX_LUT4 LUT__6034 (.I0(\useuart/r_Clock_Count[0] ), .I1(\useuart/r_Clock_Count[1] ), 
            .I2(n3960), .O(\useuart/n708 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6034.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6035 (.I0(\useuart/r_Clock_Count[0] ), .I1(\useuart/r_Clock_Count[1] ), 
            .I2(\useuart/r_Clock_Count[2] ), .I3(n3960), .O(\useuart/n711 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6035.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6036 (.I0(\useuart/r_Clock_Count[0] ), .I1(\useuart/r_Clock_Count[1] ), 
            .I2(\useuart/r_Clock_Count[2] ), .I3(\useuart/r_Clock_Count[3] ), 
            .O(n3969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__6036.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__6037 (.I0(n3969), .I1(n3960), .O(\useuart/n714 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6037.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6038 (.I0(\useuart/r_Clock_Count[0] ), .I1(\useuart/r_Clock_Count[1] ), 
            .I2(\useuart/r_Clock_Count[2] ), .I3(\useuart/r_Clock_Count[3] ), 
            .O(n3970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6038.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6039 (.I0(n3970), .I1(\useuart/r_Clock_Count[4] ), .I2(n3960), 
            .O(\useuart/n717 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6039.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6040 (.I0(n3970), .I1(\useuart/r_Clock_Count[4] ), .I2(\useuart/r_Clock_Count[5] ), 
            .I3(n3960), .O(\useuart/n720 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6040.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6041 (.I0(n3970), .I1(\useuart/r_Clock_Count[4] ), .I2(\useuart/r_Clock_Count[5] ), 
            .I3(\useuart/r_Clock_Count[6] ), .O(n3971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__6041.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__6042 (.I0(n3971), .I1(n3960), .O(\useuart/n723 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6042.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6043 (.I0(n3970), .I1(\useuart/r_Clock_Count[4] ), .I2(\useuart/r_Clock_Count[5] ), 
            .I3(\useuart/r_Clock_Count[6] ), .O(n3972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6043.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6044 (.I0(n3972), .I1(\useuart/r_Clock_Count[7] ), .I2(n3960), 
            .O(\useuart/n726 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6044.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6045 (.I0(n3972), .I1(\useuart/r_Clock_Count[7] ), .I2(\useuart/r_Clock_Count[8] ), 
            .I3(n3960), .O(\useuart/n729 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6045.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6046 (.I0(n3972), .I1(\useuart/r_Clock_Count[7] ), .I2(\useuart/r_Clock_Count[8] ), 
            .O(n3973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6046.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6047 (.I0(n3973), .I1(\useuart/r_Clock_Count[9] ), .I2(n3960), 
            .O(\useuart/n732 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6047.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6048 (.I0(n3973), .I1(\useuart/r_Clock_Count[9] ), .I2(\useuart/r_Clock_Count[10] ), 
            .I3(n3960), .O(\useuart/n735 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6048.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6049 (.I0(\useuart/r_Clock_Count[7] ), .I1(\useuart/r_Clock_Count[8] ), 
            .I2(\useuart/r_Clock_Count[9] ), .I3(\useuart/r_Clock_Count[10] ), 
            .O(n3974)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6049.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6050 (.I0(n3972), .I1(n3974), .O(n3975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6050.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6051 (.I0(n3975), .I1(\useuart/r_Clock_Count[11] ), .I2(n3960), 
            .O(\useuart/n738 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6051.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6052 (.I0(n3975), .I1(\useuart/r_Clock_Count[11] ), .I2(\useuart/r_Clock_Count[12] ), 
            .I3(n3960), .O(\useuart/n741 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6052.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6053 (.I0(\useuart/r_Bit_Index[0] ), .I1(\useuart/r_Bit_Index[1] ), 
            .I2(\useuart/r_SM_Main[1] ), .O(\useuart/n802 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6053.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6054 (.I0(\useuart/r_Bit_Index[0] ), .I1(\useuart/r_Bit_Index[1] ), 
            .I2(\useuart/r_Bit_Index[2] ), .I3(\useuart/r_SM_Main[1] ), 
            .O(\useuart/n806 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__6054.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__6055 (.I0(\useuart/LessThan_9/n26 ), .I1(\useuart/r_SM_Main[0] ), 
            .I2(\useuart/r_SM_Main[1] ), .O(\useuart/n836 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb4b4 */ ;
    defparam LUT__6055.LUTMASK = 16'hb4b4;
    EFX_LUT4 LUT__6056 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .O(n935_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__6056.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__6057 (.I0(n3881), .I1(\chunk_index[2] ), .O(n940_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__6057.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__6058 (.I0(n3881), .I1(\chunk_index[2] ), .I2(\chunk_index[3] ), 
            .O(n945_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6058.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6059 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[3] ), .O(n3976)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6059.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6060 (.I0(n3976), .I1(\chunk_index[4] ), .O(n950_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__6060.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__6061 (.I0(n3976), .I1(\chunk_index[4] ), .I2(\chunk_index[5] ), 
            .O(n955_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__6061.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__6062 (.I0(n3868), .I1(n3889), .O(n3977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6062.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6063 (.I0(n3977), .I1(\chunk_index[5] ), .I2(\state[0] ), 
            .I3(\state[1] ), .O(n868_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h88f0 */ ;
    defparam LUT__6063.LUTMASK = 16'h88f0;
    EFX_LUT4 LUT__6064 (.I0(\signature[185] ), .I1(\chunk_index[2] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n3978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b33 */ ;
    defparam LUT__6064.LUTMASK = 16'h0b33;
    EFX_LUT4 LUT__6065 (.I0(\signature[153] ), .I1(\signature[25] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n3979)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6065.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6066 (.I0(\signature[217] ), .I1(n3978), .I2(n3979), 
            .I3(\chunk_index[2] ), .O(n3980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h330d */ ;
    defparam LUT__6066.LUTMASK = 16'h330d;
    EFX_LUT4 LUT__6067 (.I0(\signature[161] ), .I1(\signature[33] ), .I2(\chunk_index[4] ), 
            .O(n3981)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6067.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6068 (.I0(\signature[225] ), .I1(\signature[97] ), .I2(\chunk_index[4] ), 
            .O(n3982)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6068.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6069 (.I0(n3982), .I1(n3981), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[2] ), .O(n3983)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6069.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6070 (.I0(n3983), .I1(n3980), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n3984)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcff5 */ ;
    defparam LUT__6070.LUTMASK = 16'hcff5;
    EFX_LUT4 LUT__6071 (.I0(\signature[145] ), .I1(\signature[129] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n3985)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6071.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6072 (.I0(n3872), .I1(n3985), .O(n3986)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6072.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6073 (.I0(\chunk_index[2] ), .I1(\chunk_index[3] ), .I2(\chunk_index[4] ), 
            .O(n3987)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6073.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6074 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .I2(\signature[57] ), 
            .I3(\chunk_index[2] ), .O(n3988)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6074.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6075 (.I0(n3987), .I1(\signature[249] ), .I2(n3988), 
            .I3(n3881), .O(n3989)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6075.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6076 (.I0(\chunk_index[0] ), .I1(\signature[113] ), .I2(\chunk_index[1] ), 
            .O(n3990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6076.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6077 (.I0(\chunk_index[0] ), .I1(\signature[209] ), .I2(\chunk_index[1] ), 
            .O(n3991)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6077.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6078 (.I0(n3991), .I1(n3870), .I2(n3858), .I3(n3990), 
            .O(n3992)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6078.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6079 (.I0(\chunk_index[2] ), .I1(\chunk_index[4] ), .I2(\chunk_index[3] ), 
            .O(n3993)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6079.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6080 (.I0(\chunk_index[0] ), .I1(\signature[81] ), .I2(\chunk_index[1] ), 
            .O(n3994)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6080.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6081 (.I0(\chunk_index[0] ), .I1(\signature[17] ), .I2(\chunk_index[1] ), 
            .O(n3995)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6081.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6082 (.I0(n3995), .I1(n3889), .I2(n3993), .I3(n3994), 
            .O(n3996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6082.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6083 (.I0(n3986), .I1(n3989), .I2(n3992), .I3(n3996), 
            .O(n3997)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6083.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6084 (.I0(\signature[201] ), .I1(\signature[169] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[3] ), .O(n3998)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6084.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6085 (.I0(\signature[105] ), .I1(\signature[9] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[3] ), .O(n3999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ff3 */ ;
    defparam LUT__6085.LUTMASK = 16'h5ff3;
    EFX_LUT4 LUT__6086 (.I0(n3999), .I1(n3998), .I2(\chunk_index[4] ), 
            .O(n4000)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6086.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6087 (.I0(\signature[1] ), .I1(\signature[137] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6087.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6088 (.I0(n3889), .I1(n3872), .I2(\chunk_index[0] ), 
            .I3(n4001), .O(n4002)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6088.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6089 (.I0(\signature[177] ), .I1(\signature[233] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4003)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6089.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6090 (.I0(n3860), .I1(n3987), .I2(n4003), .I3(\chunk_index[0] ), 
            .O(n4004)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6090.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6091 (.I0(n3874), .I1(n4000), .I2(n4002), .I3(n4004), 
            .O(n4005)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6091.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6092 (.I0(\chunk_index[4] ), .I1(\signature[121] ), .I2(n3976), 
            .O(n4006)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6092.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6093 (.I0(n3868), .I1(n3993), .I2(\signature[65] ), 
            .O(n4007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6093.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6094 (.I0(\signature[241] ), .I1(\signature[193] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[2] ), .O(n4008)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ff3 */ ;
    defparam LUT__6094.LUTMASK = 16'h5ff3;
    EFX_LUT4 LUT__6095 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .O(n4009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6095.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6096 (.I0(\chunk_index[0] ), .I1(n4008), .I2(n4009), 
            .O(n4010)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6096.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6097 (.I0(\signature[49] ), .I1(\signature[41] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4011)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6097.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6098 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .I2(\chunk_index[2] ), 
            .O(n4012)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6098.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6099 (.I0(\signature[89] ), .I1(\signature[73] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4013)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6099.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6100 (.I0(n3993), .I1(n4013), .I2(n4011), .I3(n4012), 
            .O(n4014)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__6100.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__6101 (.I0(n4006), .I1(n4007), .I2(n4010), .I3(n4014), 
            .O(n4015)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6101.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6102 (.I0(n3984), .I1(n3997), .I2(n4005), .I3(n4015), 
            .O(n827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6102.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6103 (.I0(n4012), .I1(n3874), .I2(\signature[42] ), 
            .O(n4016)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6103.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6104 (.I0(\signature[250] ), .I1(\chunk_index[2] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4017)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6104.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6105 (.I0(n3872), .I1(\signature[154] ), .I2(n4017), 
            .I3(n3881), .O(n4018)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6105.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6106 (.I0(n3889), .I1(\chunk_index[0] ), .I2(\signature[26] ), 
            .I3(\chunk_index[1] ), .O(n4019)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6106.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6107 (.I0(\signature[178] ), .I1(\signature[170] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4020)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6107.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6108 (.I0(\signature[98] ), .I1(\signature[2] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[3] ), .O(n4021)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ff3 */ ;
    defparam LUT__6108.LUTMASK = 16'h5ff3;
    EFX_LUT4 LUT__6109 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\chunk_index[4] ), 
            .O(n4022)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6109.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6110 (.I0(n4021), .I1(n4022), .I2(n4020), .I3(n3860), 
            .O(n4023)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__6110.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__6111 (.I0(n4016), .I1(n4018), .I2(n4019), .I3(n4023), 
            .O(n4024)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6111.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6112 (.I0(\chunk_index[2] ), .I1(\chunk_index[4] ), .I2(\chunk_index[3] ), 
            .I3(\signature[74] ), .O(n4025)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6112.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6113 (.I0(n3858), .I1(\signature[106] ), .I2(n4025), 
            .I3(n3874), .O(n4026)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6113.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6114 (.I0(\signature[130] ), .I1(\signature[10] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6114.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6115 (.I0(n3872), .I1(n3889), .I2(\chunk_index[0] ), 
            .I3(n4027), .O(n4028)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6115.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6116 (.I0(\signature[186] ), .I1(\signature[138] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6116.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6117 (.I0(n3872), .I1(n3860), .I2(\chunk_index[1] ), 
            .I3(n4029), .O(n4030)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6117.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6118 (.I0(\signature[146] ), .I1(\signature[58] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6118.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6119 (.I0(n3872), .I1(n4012), .I2(\chunk_index[0] ), 
            .I3(n4031), .O(n4032)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6119.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6120 (.I0(n4026), .I1(n4028), .I2(n4030), .I3(n4032), 
            .O(n4033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6120.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6121 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[34] ), 
            .O(n4034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6121.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6122 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[66] ), 
            .O(n4035)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6122.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6123 (.I0(n3993), .I1(n4035), .I2(n4012), .I3(n4034), 
            .O(n4036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6123.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6124 (.I0(\signature[210] ), .I1(\signature[162] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4037)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6124.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6125 (.I0(n3860), .I1(n3870), .I2(\chunk_index[1] ), 
            .I3(n4037), .O(n4038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6125.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6126 (.I0(\signature[82] ), .I1(\signature[218] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4039)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6126.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6127 (.I0(n3993), .I1(n3870), .I2(\chunk_index[0] ), 
            .I3(n4039), .O(n4040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6127.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6128 (.I0(\signature[202] ), .I1(\signature[122] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4041)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6128.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6129 (.I0(n3870), .I1(n3858), .I2(\chunk_index[1] ), 
            .I3(n4041), .O(n4042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6129.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6130 (.I0(n4038), .I1(n4040), .I2(n4042), .I3(n4036), 
            .O(n4043)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6130.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6131 (.I0(\signature[242] ), .I1(\signature[234] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6131.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6132 (.I0(n4044), .I1(n3987), .O(n4045)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6132.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6133 (.I0(\chunk_index[2] ), .I1(\signature[194] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6133.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6134 (.I0(\chunk_index[0] ), .I1(\signature[18] ), .I2(\chunk_index[1] ), 
            .O(n4047)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6134.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6135 (.I0(n4047), .I1(n3889), .I2(n3868), .I3(n4046), 
            .O(n4048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6135.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6136 (.I0(\signature[114] ), .I1(\signature[90] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4049)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6136.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6137 (.I0(n3858), .I1(n3993), .I2(\chunk_index[0] ), 
            .I3(n4049), .O(n4050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6137.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6138 (.I0(\signature[226] ), .I1(\signature[50] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4051)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6138.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6139 (.I0(n3987), .I1(n4012), .I2(\chunk_index[1] ), 
            .I3(n4051), .O(n4052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6139.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6140 (.I0(n4045), .I1(n4050), .I2(n4052), .I3(n4048), 
            .O(n4053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6140.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6141 (.I0(n4024), .I1(n4033), .I2(n4043), .I3(n4053), 
            .O(n826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6141.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6142 (.I0(n3860), .I1(\signature[179] ), .I2(\signature[19] ), 
            .I3(n3889), .O(n4054)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6142.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6143 (.I0(n3872), .I1(n3881), .I2(\signature[155] ), 
            .O(n4055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6143.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6144 (.I0(\signature[251] ), .I1(\chunk_index[2] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4056)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6144.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6145 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .I2(\signature[51] ), 
            .I3(\chunk_index[2] ), .O(n4057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6145.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6146 (.I0(n4057), .I1(n4056), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4058)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6146.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6147 (.I0(n3877), .I1(n4054), .I2(n4055), .I3(n4058), 
            .O(n4059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__6147.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__6148 (.I0(\signature[243] ), .I1(\signature[235] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6148.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6149 (.I0(n3868), .I1(\signature[227] ), .I2(n4060), 
            .I3(n3987), .O(n4061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__6149.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__6150 (.I0(\signature[59] ), .I1(\signature[43] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4062)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6150.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6151 (.I0(n3868), .I1(\signature[35] ), .I2(n4062), 
            .I3(n4012), .O(n4063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6151.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6152 (.I0(\chunk_index[4] ), .I1(\chunk_index[2] ), .I2(\chunk_index[3] ), 
            .I3(\signature[123] ), .O(n4064)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6152.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6153 (.I0(n3860), .I1(\signature[187] ), .I2(n4064), 
            .I3(n3881), .O(n4065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6153.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6154 (.I0(\chunk_index[3] ), .I1(\chunk_index[2] ), .I2(\signature[163] ), 
            .I3(\chunk_index[4] ), .O(n4066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6154.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6155 (.I0(\signature[195] ), .I1(\signature[99] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[4] ), .O(n4067)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6155.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6156 (.I0(n4067), .I1(n3892), .I2(n3868), .I3(n4066), 
            .O(n4068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__6156.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__6157 (.I0(n4061), .I1(n4063), .I2(n4065), .I3(n4068), 
            .O(n4069)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6157.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6158 (.I0(\signature[83] ), .I1(\signature[91] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6158.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6159 (.I0(\signature[27] ), .I1(\signature[11] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6159.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6160 (.I0(n4071), .I1(n3889), .I2(n3993), .I3(n4070), 
            .O(n4072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6160.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6161 (.I0(n3868), .I1(n3993), .I2(\signature[67] ), 
            .O(n4073)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6161.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6162 (.I0(\signature[115] ), .I1(\signature[107] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6162.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6163 (.I0(\signature[147] ), .I1(\signature[139] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6163.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6164 (.I0(n4075), .I1(n3872), .I2(n4074), .I3(n3858), 
            .O(n4076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__6164.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__6165 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[3] ), 
            .O(n4077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6165.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6166 (.I0(\signature[211] ), .I1(\signature[219] ), .I2(\chunk_index[0] ), 
            .O(n4078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6166.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6167 (.I0(\chunk_index[2] ), .I1(\chunk_index[1] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4079)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6167.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6168 (.I0(n4078), .I1(n4079), .I2(n3889), .I3(n4077), 
            .O(n4080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__6168.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__6169 (.I0(n4073), .I1(n4072), .I2(n4076), .I3(n4080), 
            .O(n4081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6169.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6170 (.I0(n3870), .I1(\signature[203] ), .I2(\signature[75] ), 
            .I3(n3993), .O(n4082)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6170.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6171 (.I0(\signature[131] ), .I1(\signature[171] ), .I2(\chunk_index[0] ), 
            .O(n4083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6171.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6172 (.I0(n3872), .I1(n3860), .I2(n4083), .I3(\chunk_index[0] ), 
            .O(n4084)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6172.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6173 (.I0(\chunk_index[1] ), .I1(n4084), .I2(n4082), 
            .I3(n3874), .O(n4085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__6173.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__6174 (.I0(n4059), .I1(n4069), .I2(n4081), .I3(n4085), 
            .O(n825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6174.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6175 (.I0(\signature[220] ), .I1(\signature[92] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6175.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6176 (.I0(\signature[156] ), .I1(\signature[188] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[2] ), .O(n4087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf305 */ ;
    defparam LUT__6176.LUTMASK = 16'hf305;
    EFX_LUT4 LUT__6177 (.I0(n4086), .I1(n4087), .O(n4088)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6177.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6178 (.I0(\signature[204] ), .I1(\signature[140] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[3] ), .O(n4089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__6178.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__6179 (.I0(\chunk_index[2] ), .I1(\signature[236] ), .I2(n4089), 
            .I3(\chunk_index[4] ), .O(n4090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6179.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6180 (.I0(n4090), .I1(n4088), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6180.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6181 (.I0(\signature[84] ), .I1(\signature[76] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6181.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6182 (.I0(n4092), .I1(n3993), .O(n4093)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6182.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6183 (.I0(\chunk_index[0] ), .I1(\signature[52] ), .I2(\chunk_index[1] ), 
            .O(n4094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6183.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6184 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[228] ), 
            .I3(\chunk_index[2] ), .O(n4095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6184.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6185 (.I0(n4094), .I1(n4012), .I2(n4009), .I3(n4095), 
            .O(n4096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6185.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6186 (.I0(\signature[116] ), .I1(\signature[100] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4097)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6186.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6187 (.I0(n3874), .I1(\signature[108] ), .I2(n4097), 
            .I3(n3858), .O(n4098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6187.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6188 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[2] ), .O(n4099)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6188.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6189 (.I0(\signature[164] ), .I1(\signature[36] ), .I2(\chunk_index[4] ), 
            .I3(n4099), .O(n4100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6189.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6190 (.I0(n4093), .I1(n4098), .I2(n4100), .I3(n4096), 
            .O(n4101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6190.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6191 (.I0(\signature[180] ), .I1(\signature[172] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6191.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6192 (.I0(n4102), .I1(n3860), .O(n4103)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6192.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6193 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[132] ), 
            .O(n4104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6193.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6194 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[4] ), 
            .O(n4105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6194.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6195 (.I0(n3889), .I1(n4105), .I2(n3872), .I3(n4104), 
            .O(n4106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6195.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6196 (.I0(\signature[20] ), .I1(\signature[44] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4107)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6196.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6197 (.I0(n3889), .I1(n4012), .I2(n4107), .I3(\chunk_index[0] ), 
            .O(n4108)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6197.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6198 (.I0(\signature[196] ), .I1(\signature[124] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4109)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff5 */ ;
    defparam LUT__6198.LUTMASK = 16'h3ff5;
    EFX_LUT4 LUT__6199 (.I0(n3870), .I1(n3858), .I2(n4109), .I3(\chunk_index[0] ), 
            .O(n4110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6199.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6200 (.I0(n4103), .I1(n4108), .I2(n4110), .I3(n4106), 
            .O(n4111)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6200.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6201 (.I0(\signature[28] ), .I1(\signature[12] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4112)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6201.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6202 (.I0(n3889), .I1(n4112), .O(n4113)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6202.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6203 (.I0(\signature[244] ), .I1(\signature[212] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[1] ), .O(n4114)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6203.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6204 (.I0(\chunk_index[0] ), .I1(n4114), .I2(n4009), 
            .O(n4115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6204.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6205 (.I0(\signature[68] ), .I1(\signature[60] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4116)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff5 */ ;
    defparam LUT__6205.LUTMASK = 16'h3ff5;
    EFX_LUT4 LUT__6206 (.I0(n3993), .I1(n4012), .I2(n4116), .I3(\chunk_index[0] ), 
            .O(n4117)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6206.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6207 (.I0(\signature[148] ), .I1(\signature[252] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6207.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6208 (.I0(n3872), .I1(n3987), .I2(\chunk_index[0] ), 
            .I3(n4118), .O(n4119)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6208.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6209 (.I0(n4113), .I1(n4115), .I2(n4117), .I3(n4119), 
            .O(n4120)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6209.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6210 (.I0(n4091), .I1(n4101), .I2(n4111), .I3(n4120), 
            .O(n824)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6210.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6211 (.I0(\chunk_index[2] ), .I1(\signature[205] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6211.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6212 (.I0(\signature[141] ), .I1(n3872), .I2(n4121), 
            .I3(n3874), .O(n4122)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6212.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6213 (.I0(\signature[229] ), .I1(\signature[213] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[2] ), .O(n4123)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6213.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6214 (.I0(n4123), .I1(\chunk_index[3] ), .I2(\chunk_index[4] ), 
            .I3(\chunk_index[0] ), .O(n4124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__6214.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__6215 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .I2(\signature[61] ), 
            .I3(\chunk_index[2] ), .O(n4125)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6215.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6216 (.I0(\signature[189] ), .I1(n3860), .I2(n4125), 
            .I3(n3881), .O(n4126)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6216.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6217 (.I0(n4122), .I1(n4124), .I2(n4126), .O(n4127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6217.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6218 (.I0(\chunk_index[2] ), .I1(\chunk_index[3] ), .I2(\signature[133] ), 
            .I3(\chunk_index[4] ), .O(n4128)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6218.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6219 (.I0(n4012), .I1(\signature[53] ), .I2(n4128), 
            .I3(\chunk_index[1] ), .O(n4129)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__6219.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__6220 (.I0(\signature[253] ), .I1(\signature[125] ), .I2(\chunk_index[4] ), 
            .I3(n3976), .O(n4130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6220.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6221 (.I0(n3868), .I1(n3889), .I2(\signature[5] ), .O(n4131)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6221.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6222 (.I0(\chunk_index[0] ), .I1(n4129), .I2(n4130), 
            .I3(n4131), .O(n4132)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__6222.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__6223 (.I0(\signature[197] ), .I1(\signature[45] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6223.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6224 (.I0(n3870), .I1(n4012), .I2(\chunk_index[0] ), 
            .I3(n4133), .O(n4134)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6224.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6225 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[69] ), 
            .O(n4135)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6225.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6226 (.I0(\signature[101] ), .I1(\signature[109] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6226.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6227 (.I0(n4135), .I1(n3993), .I2(n3858), .I3(n4136), 
            .O(n4137)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6227.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6228 (.I0(\signature[93] ), .I1(\signature[77] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h503f */ ;
    defparam LUT__6228.LUTMASK = 16'h503f;
    EFX_LUT4 LUT__6229 (.I0(\signature[85] ), .I1(\chunk_index[0] ), .I2(n4138), 
            .I3(n3993), .O(n4139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__6229.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__6230 (.I0(\signature[181] ), .I1(\signature[173] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6230.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6231 (.I0(\signature[245] ), .I1(\signature[237] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6231.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6232 (.I0(n4141), .I1(n3987), .I2(n4140), .I3(n3860), 
            .O(n4142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__6232.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__6233 (.I0(n4134), .I1(n4139), .I2(n4137), .I3(n4142), 
            .O(n4143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6233.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6234 (.I0(\chunk_index[3] ), .I1(\chunk_index[4] ), .I2(\signature[37] ), 
            .I3(\chunk_index[2] ), .O(n4144)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6234.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6235 (.I0(n3860), .I1(\signature[165] ), .I2(n4144), 
            .I3(n3868), .O(n4145)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6235.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6236 (.I0(\signature[13] ), .I1(\signature[21] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0 */ ;
    defparam LUT__6236.LUTMASK = 16'hfac0;
    EFX_LUT4 LUT__6237 (.I0(\signature[29] ), .I1(n3881), .I2(n4146), 
            .I3(n3889), .O(n4147)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6237.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6238 (.I0(\chunk_index[2] ), .I1(\chunk_index[3] ), .I2(\signature[149] ), 
            .I3(\chunk_index[4] ), .O(n4148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6238.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6239 (.I0(n3858), .I1(\signature[117] ), .I2(n4148), 
            .I3(n3877), .O(n4149)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6239.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6240 (.I0(\chunk_index[2] ), .I1(\signature[221] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6240.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6241 (.I0(n3872), .I1(\signature[157] ), .I2(n4150), 
            .I3(n3881), .O(n4151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6241.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6242 (.I0(n4145), .I1(n4147), .I2(n4149), .I3(n4151), 
            .O(n4152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6242.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6243 (.I0(n4127), .I1(n4132), .I2(n4143), .I3(n4152), 
            .O(n823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6243.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6244 (.I0(\signature[38] ), .I1(\signature[6] ), .I2(\chunk_index[4] ), 
            .I3(\chunk_index[2] ), .O(n4153)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h05f3 */ ;
    defparam LUT__6244.LUTMASK = 16'h05f3;
    EFX_LUT4 LUT__6245 (.I0(\signature[166] ), .I1(\signature[230] ), .I2(\chunk_index[4] ), 
            .I3(\chunk_index[3] ), .O(n4154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3f50 */ ;
    defparam LUT__6245.LUTMASK = 16'h3f50;
    EFX_LUT4 LUT__6246 (.I0(\signature[102] ), .I1(\signature[126] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4155)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff5 */ ;
    defparam LUT__6246.LUTMASK = 16'h3ff5;
    EFX_LUT4 LUT__6247 (.I0(n3877), .I1(\signature[118] ), .I2(n4155), 
            .I3(n3858), .O(n4156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__6247.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__6248 (.I0(n4154), .I1(n4153), .I2(n3868), .I3(n4156), 
            .O(n4157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6248.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6249 (.I0(n3877), .I1(n3889), .I2(\signature[22] ), 
            .O(n4158)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6249.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6250 (.I0(\signature[150] ), .I1(\signature[142] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6250.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6251 (.I0(n3868), .I1(\signature[134] ), .I2(n4159), 
            .I3(n3872), .O(n4160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__6251.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__6252 (.I0(\signature[254] ), .I1(\signature[238] ), .I2(\chunk_index[1] ), 
            .O(n4161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6252.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6253 (.I0(\signature[86] ), .I1(\signature[78] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6253.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6254 (.I0(n4162), .I1(n3993), .I2(n4161), .I3(n3897), 
            .O(n4163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__6254.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__6255 (.I0(\signature[214] ), .I1(\signature[70] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6255.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6256 (.I0(n3993), .I1(n3870), .I2(\chunk_index[1] ), 
            .I3(n4164), .O(n4165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6256.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6257 (.I0(n4158), .I1(n4160), .I2(n4165), .I3(n4163), 
            .O(n4166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6257.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6258 (.I0(\signature[246] ), .I1(\signature[222] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[2] ), .O(n4167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6258.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6259 (.I0(n4167), .I1(n4009), .I2(\chunk_index[1] ), 
            .O(n4168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6259.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6260 (.I0(\signature[54] ), .I1(\signature[174] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6260.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6261 (.I0(n4012), .I1(n3860), .I2(n4169), .I3(\chunk_index[0] ), 
            .O(n4170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6261.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6262 (.I0(\signature[110] ), .I1(\signature[62] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6262.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6263 (.I0(n3858), .I1(n4012), .I2(\chunk_index[1] ), 
            .I3(n4171), .O(n4172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6263.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6264 (.I0(\signature[190] ), .I1(\signature[46] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6264.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6265 (.I0(n4012), .I1(n3860), .I2(\chunk_index[1] ), 
            .I3(n4173), .O(n4174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6265.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6266 (.I0(n4168), .I1(n4170), .I2(n4172), .I3(n4174), 
            .O(n4175)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6266.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6267 (.I0(\signature[30] ), .I1(\signature[14] ), .I2(\chunk_index[1] ), 
            .O(n4176)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6267.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6268 (.I0(\chunk_index[1] ), .I1(\chunk_index[2] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6268.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6269 (.I0(n4177), .I1(\signature[206] ), .I2(n4176), 
            .I3(n3889), .O(n4178)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__6269.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__6270 (.I0(\signature[198] ), .I1(\signature[158] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4179)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff5 */ ;
    defparam LUT__6270.LUTMASK = 16'h3ff5;
    EFX_LUT4 LUT__6271 (.I0(n3870), .I1(n3872), .I2(n4179), .I3(\chunk_index[0] ), 
            .O(n4180)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6271.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6272 (.I0(\signature[182] ), .I1(\signature[94] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4181)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6272.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6273 (.I0(n3860), .I1(n3993), .I2(\chunk_index[0] ), 
            .I3(n4181), .O(n4182)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6273.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6274 (.I0(\chunk_index[0] ), .I1(n4178), .I2(n4180), 
            .I3(n4182), .O(n4183)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__6274.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__6275 (.I0(n4157), .I1(n4166), .I2(n4175), .I3(n4183), 
            .O(n822)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6275.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6276 (.I0(\signature[71] ), .I1(n3993), .I2(n3860), 
            .I3(\signature[167] ), .O(n4184)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6276.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6277 (.I0(\signature[55] ), .I1(\signature[47] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4185)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6277.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6278 (.I0(\signature[39] ), .I1(\signature[63] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4186)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ff5 */ ;
    defparam LUT__6278.LUTMASK = 16'h3ff5;
    EFX_LUT4 LUT__6279 (.I0(n4186), .I1(n4185), .I2(n4012), .O(n4187)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__6279.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__6280 (.I0(\signature[119] ), .I1(\signature[111] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4188)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6280.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6281 (.I0(\chunk_index[0] ), .I1(\signature[215] ), .I2(\chunk_index[1] ), 
            .O(n4189)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6281.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6282 (.I0(n4189), .I1(n3870), .I2(n4188), .I3(n3858), 
            .O(n4190)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__6282.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__6283 (.I0(n3868), .I1(n4184), .I2(n4187), .I3(n4190), 
            .O(n4191)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6283.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6284 (.I0(\signature[255] ), .I1(\signature[127] ), .I2(\chunk_index[4] ), 
            .I3(n3976), .O(n4192)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6284.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6285 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[103] ), 
            .O(n4193)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6285.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6286 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[135] ), 
            .O(n4194)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6286.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6287 (.I0(n4194), .I1(n3872), .I2(n3858), .I3(n4193), 
            .O(n4195)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6287.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6288 (.I0(\signature[151] ), .I1(\signature[7] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4196)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6288.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6289 (.I0(n3889), .I1(n3872), .I2(\chunk_index[1] ), 
            .I3(n4196), .O(n4197)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6289.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6290 (.I0(\signature[87] ), .I1(\signature[95] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4198)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6290.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6291 (.I0(\chunk_index[0] ), .I1(\chunk_index[1] ), .I2(\signature[199] ), 
            .O(n4199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6291.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6292 (.I0(n4199), .I1(n3870), .I2(n3993), .I3(n4198), 
            .O(n4200)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6292.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6293 (.I0(n4192), .I1(n4197), .I2(n4195), .I3(n4200), 
            .O(n4201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6293.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6294 (.I0(n3889), .I1(n3874), .I2(\signature[15] ), 
            .O(n4202)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6294.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6295 (.I0(n3860), .I1(n3877), .I2(\signature[183] ), 
            .O(n4203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6295.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6296 (.I0(\signature[239] ), .I1(\signature[223] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[2] ), .O(n4204)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6296.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6297 (.I0(n4204), .I1(\chunk_index[0] ), .I2(\chunk_index[3] ), 
            .I3(\chunk_index[4] ), .O(n4205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6297.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6298 (.I0(\chunk_index[2] ), .I1(\chunk_index[3] ), .I2(\chunk_index[4] ), 
            .I3(\signature[23] ), .O(n4206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6298.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6299 (.I0(\chunk_index[3] ), .I1(\chunk_index[2] ), .I2(\signature[191] ), 
            .I3(\chunk_index[4] ), .O(n4207)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6299.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6300 (.I0(n4207), .I1(n4206), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6300.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6301 (.I0(n4202), .I1(n4203), .I2(n4205), .I3(n4208), 
            .O(n4209)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6301.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6302 (.I0(\signature[79] ), .I1(\signature[31] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[3] ), .O(n4210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6302.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6303 (.I0(n4210), .I1(\chunk_index[2] ), .I2(\chunk_index[4] ), 
            .I3(\chunk_index[0] ), .O(n4211)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6303.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6304 (.I0(\signature[231] ), .I1(\signature[175] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[3] ), .O(n4212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6304.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6305 (.I0(n4212), .I1(\chunk_index[1] ), .I2(\chunk_index[2] ), 
            .I3(\chunk_index[4] ), .O(n4213)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6305.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6306 (.I0(\signature[247] ), .I1(\signature[143] ), .I2(\chunk_index[0] ), 
            .I3(\chunk_index[1] ), .O(n4214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf53f */ ;
    defparam LUT__6306.LUTMASK = 16'hf53f;
    EFX_LUT4 LUT__6307 (.I0(n3987), .I1(n3872), .I2(n4214), .I3(\chunk_index[0] ), 
            .O(n4215)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6307.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6308 (.I0(\signature[207] ), .I1(\signature[159] ), .I2(\chunk_index[1] ), 
            .I3(\chunk_index[0] ), .O(n4216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6308.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6309 (.I0(n3870), .I1(n3872), .I2(\chunk_index[1] ), 
            .I3(n4216), .O(n4217)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6309.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6310 (.I0(n4211), .I1(n4213), .I2(n4215), .I3(n4217), 
            .O(n4218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6310.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6311 (.I0(n4191), .I1(n4201), .I2(n4209), .I3(n4218), 
            .O(n821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6311.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6312 (.I0(\useone/a[1] ), .I1(\useone/a[12] ), .I2(\useone/a[21] ), 
            .O(n3421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6312.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6313 (.I0(\useone/a[31] ), .I1(\useone/b[31] ), .I2(\useone/c[31] ), 
            .O(n3422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__6313.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__6314 (.I0(\useone/a[0] ), .I1(\useone/a[11] ), .I2(\useone/a[20] ), 
            .O(n3424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6314.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6315 (.I0(\useone/a[30] ), .I1(\useone/b[30] ), .I2(\useone/c[30] ), 
            .O(n3425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd4d4 */ ;
    defparam LUT__6315.LUTMASK = 16'hd4d4;
    EFX_LUT4 LUT__6316 (.I0(\useone/a[10] ), .I1(\useone/a[19] ), .I2(\useone/a[31] ), 
            .O(n3427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6316.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6317 (.I0(\useone/a[29] ), .I1(\useone/b[29] ), .I2(\useone/c[29] ), 
            .O(n3428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1717 */ ;
    defparam LUT__6317.LUTMASK = 16'h1717;
    EFX_LUT4 LUT__6318 (.I0(\useone/a[9] ), .I1(\useone/a[18] ), .I2(\useone/a[30] ), 
            .O(n3430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6318.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6319 (.I0(\useone/a[28] ), .I1(\useone/b[28] ), .I2(\useone/c[28] ), 
            .O(n3431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__6319.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__6320 (.I0(\useone/a[8] ), .I1(\useone/a[17] ), .I2(\useone/a[29] ), 
            .O(n3433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6320.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6321 (.I0(\useone/a[27] ), .I1(\useone/b[27] ), .I2(\useone/c[27] ), 
            .O(n3434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1717 */ ;
    defparam LUT__6321.LUTMASK = 16'h1717;
    EFX_LUT4 LUT__6322 (.I0(\useone/a[7] ), .I1(\useone/a[16] ), .I2(\useone/a[28] ), 
            .O(n3436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6322.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6323 (.I0(\useone/a[26] ), .I1(\useone/c[26] ), .I2(\useone/b[26] ), 
            .O(n3437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__6323.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__6324 (.I0(\useone/a[6] ), .I1(\useone/a[15] ), .I2(\useone/a[27] ), 
            .O(n3439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6324.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6325 (.I0(\useone/a[25] ), .I1(\useone/b[25] ), .I2(\useone/c[25] ), 
            .O(n3440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6325.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6326 (.I0(\useone/a[5] ), .I1(\useone/a[14] ), .I2(\useone/a[26] ), 
            .O(n3442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6326.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6327 (.I0(\useone/a[24] ), .I1(\useone/b[24] ), .I2(\useone/c[24] ), 
            .O(n3443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__6327.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__6328 (.I0(\useone/a[4] ), .I1(\useone/a[13] ), .I2(\useone/a[25] ), 
            .O(n3445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6328.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6329 (.I0(\useone/a[23] ), .I1(\useone/b[23] ), .I2(\useone/c[23] ), 
            .O(n3446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8e8 */ ;
    defparam LUT__6329.LUTMASK = 16'he8e8;
    EFX_LUT4 LUT__6330 (.I0(\useone/a[3] ), .I1(\useone/a[12] ), .I2(\useone/a[24] ), 
            .O(n3448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6330.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6331 (.I0(\useone/a[22] ), .I1(\useone/b[22] ), .I2(\useone/c[22] ), 
            .O(n3449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__6331.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__6332 (.I0(\useone/a[2] ), .I1(\useone/a[11] ), .I2(\useone/a[23] ), 
            .O(n3451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6332.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6333 (.I0(\useone/a[21] ), .I1(\useone/b[21] ), .I2(\useone/c[21] ), 
            .O(n3452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__6333.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__6334 (.I0(\useone/a[1] ), .I1(\useone/a[10] ), .I2(\useone/a[22] ), 
            .O(n3454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6334.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6335 (.I0(\useone/a[20] ), .I1(\useone/b[20] ), .I2(\useone/c[20] ), 
            .O(n3455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8e8 */ ;
    defparam LUT__6335.LUTMASK = 16'he8e8;
    EFX_LUT4 LUT__6336 (.I0(\useone/a[0] ), .I1(\useone/a[9] ), .I2(\useone/a[21] ), 
            .O(n3457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6336.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6337 (.I0(\useone/a[19] ), .I1(\useone/c[19] ), .I2(\useone/b[19] ), 
            .O(n3458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6337.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6338 (.I0(\useone/a[8] ), .I1(\useone/a[20] ), .I2(\useone/a[31] ), 
            .O(n3460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6338.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6339 (.I0(\useone/a[18] ), .I1(\useone/b[18] ), .I2(\useone/c[18] ), 
            .O(n3461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__6339.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__6340 (.I0(\useone/a[7] ), .I1(\useone/a[19] ), .I2(\useone/a[30] ), 
            .O(n3463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6340.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6341 (.I0(\useone/a[17] ), .I1(\useone/b[17] ), .I2(\useone/c[17] ), 
            .O(n3464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__6341.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__6342 (.I0(\useone/a[6] ), .I1(\useone/a[18] ), .I2(\useone/a[29] ), 
            .O(n3466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6342.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6343 (.I0(\useone/a[16] ), .I1(\useone/b[16] ), .I2(\useone/c[16] ), 
            .O(n3467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6343.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6344 (.I0(\useone/a[5] ), .I1(\useone/a[17] ), .I2(\useone/a[28] ), 
            .O(n3469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6344.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6345 (.I0(\useone/a[15] ), .I1(\useone/b[15] ), .I2(\useone/c[15] ), 
            .O(n3470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1717 */ ;
    defparam LUT__6345.LUTMASK = 16'h1717;
    EFX_LUT4 LUT__6346 (.I0(\useone/a[4] ), .I1(\useone/a[16] ), .I2(\useone/a[27] ), 
            .O(n3472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6346.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6347 (.I0(\useone/a[14] ), .I1(\useone/c[14] ), .I2(\useone/b[14] ), 
            .O(n3473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6347.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6348 (.I0(\useone/a[3] ), .I1(\useone/a[15] ), .I2(\useone/a[26] ), 
            .O(n3475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6348.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6349 (.I0(\useone/a[13] ), .I1(\useone/b[13] ), .I2(\useone/c[13] ), 
            .O(n3476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1717 */ ;
    defparam LUT__6349.LUTMASK = 16'h1717;
    EFX_LUT4 LUT__6350 (.I0(\useone/a[2] ), .I1(\useone/a[14] ), .I2(\useone/a[25] ), 
            .O(n3478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6350.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6351 (.I0(\useone/a[12] ), .I1(\useone/c[12] ), .I2(\useone/b[12] ), 
            .O(n3479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__6351.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__6352 (.I0(\useone/a[1] ), .I1(\useone/a[13] ), .I2(\useone/a[24] ), 
            .O(n3481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6352.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6353 (.I0(\useone/a[11] ), .I1(\useone/b[11] ), .I2(\useone/c[11] ), 
            .O(n3482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__6353.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__6354 (.I0(\useone/a[0] ), .I1(\useone/a[12] ), .I2(\useone/a[23] ), 
            .O(n3484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6354.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6355 (.I0(\useone/a[10] ), .I1(\useone/b[10] ), .I2(\useone/c[10] ), 
            .O(n3485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6355.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6356 (.I0(\useone/a[11] ), .I1(\useone/a[22] ), .I2(\useone/a[31] ), 
            .O(n3487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6356.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6357 (.I0(\useone/a[9] ), .I1(\useone/b[9] ), .I2(\useone/c[9] ), 
            .O(n3488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1717 */ ;
    defparam LUT__6357.LUTMASK = 16'h1717;
    EFX_LUT4 LUT__6358 (.I0(\useone/a[10] ), .I1(\useone/a[21] ), .I2(\useone/a[30] ), 
            .O(n3490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6358.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6359 (.I0(\useone/a[8] ), .I1(\useone/c[8] ), .I2(\useone/b[8] ), 
            .O(n3491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__6359.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__6360 (.I0(\useone/a[9] ), .I1(\useone/a[20] ), .I2(\useone/a[29] ), 
            .O(n3493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6360.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6361 (.I0(\useone/a[7] ), .I1(\useone/b[7] ), .I2(\useone/c[7] ), 
            .O(n3494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__6361.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__6362 (.I0(\useone/a[8] ), .I1(\useone/a[19] ), .I2(\useone/a[28] ), 
            .O(n3496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6362.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6363 (.I0(\useone/a[6] ), .I1(\useone/c[6] ), .I2(\useone/b[6] ), 
            .O(n3497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6363.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6364 (.I0(\useone/a[7] ), .I1(\useone/a[18] ), .I2(\useone/a[27] ), 
            .O(n3499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6364.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6365 (.I0(\useone/a[5] ), .I1(\useone/c[5] ), .I2(\useone/b[5] ), 
            .O(n3500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6365.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6366 (.I0(\useone/a[6] ), .I1(\useone/a[17] ), .I2(\useone/a[26] ), 
            .O(n3502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6366.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6367 (.I0(\useone/a[4] ), .I1(\useone/c[4] ), .I2(\useone/b[4] ), 
            .O(n3503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb2b2 */ ;
    defparam LUT__6367.LUTMASK = 16'hb2b2;
    EFX_LUT4 LUT__6368 (.I0(\useone/a[5] ), .I1(\useone/a[16] ), .I2(\useone/a[25] ), 
            .O(n3505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6368.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6369 (.I0(\useone/a[3] ), .I1(\useone/b[3] ), .I2(\useone/c[3] ), 
            .O(n3506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he8e8 */ ;
    defparam LUT__6369.LUTMASK = 16'he8e8;
    EFX_LUT4 LUT__6370 (.I0(\useone/a[4] ), .I1(\useone/a[15] ), .I2(\useone/a[24] ), 
            .O(n3508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6370.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6371 (.I0(\useone/a[2] ), .I1(\useone/b[2] ), .I2(\useone/c[2] ), 
            .O(n3509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6371.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6372 (.I0(\useone/a[3] ), .I1(\useone/a[14] ), .I2(\useone/a[23] ), 
            .O(n3511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6372.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6373 (.I0(\useone/a[1] ), .I1(\useone/c[1] ), .I2(\useone/b[1] ), 
            .O(n3512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7171 */ ;
    defparam LUT__6373.LUTMASK = 16'h7171;
    EFX_LUT4 LUT__6374 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[2] ), .O(n4219)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8e53 */ ;
    defparam LUT__6374.LUTMASK = 16'h8e53;
    EFX_LUT4 LUT__6375 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[4] ), 
            .O(n4220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6375.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6376 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .O(n4221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6376.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6377 (.I0(n4221), .I1(n4220), .I2(n3914), .O(n4222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6377.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6378 (.I0(\useone/round_flag[1] ), .I1(n4219), .I2(n4222), 
            .O(n4223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6378.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6379 (.I0(n1191_2), .I1(\useone/round_flag[5] ), .O(n4224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6379.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6380 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[2] ), .O(n4225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbdc3 */ ;
    defparam LUT__6380.LUTMASK = 16'hbdc3;
    EFX_LUT4 LUT__6381 (.I0(\useone/round_flag[5] ), .I1(\useone/round_flag[4] ), 
            .O(n4226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6381.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6382 (.I0(n4226), .I1(n1191_2), .O(n4227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6382.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6383 (.I0(n4225), .I1(n4227), .I2(n4223), .I3(n4224), 
            .O(n3515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf444 */ ;
    defparam LUT__6383.LUTMASK = 16'hf444;
    EFX_LUT4 LUT__6384 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[1] ), 
            .O(n4228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6384.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6385 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[3] ), .O(n4229)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6385.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6386 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[4] ), .O(n4230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcda3 */ ;
    defparam LUT__6386.LUTMASK = 16'hcda3;
    EFX_LUT4 LUT__6387 (.I0(n4229), .I1(n4228), .I2(n4230), .I3(\useone/round_flag[0] ), 
            .O(n4231)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6387.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6388 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(n4231), .O(n4232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__6388.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__6389 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4233)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3ec */ ;
    defparam LUT__6389.LUTMASK = 16'hc3ec;
    EFX_LUT4 LUT__6390 (.I0(n3909), .I1(\useone/round_flag[4] ), .I2(n4233), 
            .I3(\useone/round_flag[2] ), .O(n4234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__6390.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__6391 (.I0(n4234), .I1(n4232), .I2(\useone/round_flag[5] ), 
            .I3(n1191_2), .O(n3518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6391.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6392 (.I0(\useone/round_flag[0] ), .I1(n3910), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[4] ), .O(n4235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7af3 */ ;
    defparam LUT__6392.LUTMASK = 16'h7af3;
    EFX_LUT4 LUT__6393 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[4] ), .O(n4236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1401 */ ;
    defparam LUT__6393.LUTMASK = 16'h1401;
    EFX_LUT4 LUT__6394 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[0] ), .O(n4237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hec0b */ ;
    defparam LUT__6394.LUTMASK = 16'hec0b;
    EFX_LUT4 LUT__6395 (.I0(n4236), .I1(\useone/round_flag[2] ), .I2(n4237), 
            .O(n4238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3d3d */ ;
    defparam LUT__6395.LUTMASK = 16'h3d3d;
    EFX_LUT4 LUT__6396 (.I0(n3931), .I1(\useone/round_flag[4] ), .I2(n4224), 
            .I3(n4238), .O(n4239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd000 */ ;
    defparam LUT__6396.LUTMASK = 16'hd000;
    EFX_LUT4 LUT__6397 (.I0(\useone/round_flag[5] ), .I1(n1191_2), .O(n4240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6397.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6398 (.I0(n4236), .I1(n4235), .I2(n4240), .I3(n4239), 
            .O(n3521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__6398.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__6399 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[3] ), .O(n4241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcab2 */ ;
    defparam LUT__6399.LUTMASK = 16'hcab2;
    EFX_LUT4 LUT__6400 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[1] ), .O(n4242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6400.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6401 (.I0(n4242), .I1(n4241), .I2(\useone/round_flag[4] ), 
            .O(n4243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6401.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6402 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[1] ), .O(n4244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4fba */ ;
    defparam LUT__6402.LUTMASK = 16'h4fba;
    EFX_LUT4 LUT__6403 (.I0(\useone/round_flag[2] ), .I1(n3928), .I2(n4228), 
            .I3(\useone/round_flag[4] ), .O(n4245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6403.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6404 (.I0(\useone/round_flag[4] ), .I1(n4244), .I2(n4245), 
            .I3(\useone/round_flag[5] ), .O(n4246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__6404.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__6405 (.I0(\useone/round_flag[5] ), .I1(n4243), .I2(n4246), 
            .I3(n1191_2), .O(n3524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__6405.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__6406 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc4fc */ ;
    defparam LUT__6406.LUTMASK = 16'hc4fc;
    EFX_LUT4 LUT__6407 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .O(n4248)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6407.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6408 (.I0(\useone/round_flag[2] ), .I1(n4248), .I2(\useone/round_flag[0] ), 
            .I3(\useone/round_flag[4] ), .O(n4249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c05 */ ;
    defparam LUT__6408.LUTMASK = 16'h0c05;
    EFX_LUT4 LUT__6409 (.I0(n4247), .I1(\useone/round_flag[3] ), .I2(n4249), 
            .O(n4250)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__6409.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6410 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[2] ), .O(n4251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8e53 */ ;
    defparam LUT__6410.LUTMASK = 16'h8e53;
    EFX_LUT4 LUT__6411 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[4] ), 
            .O(n4252)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6411.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6412 (.I0(n3910), .I1(n4252), .I2(n4251), .I3(\useone/round_flag[4] ), 
            .O(n4253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__6412.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__6413 (.I0(n4253), .I1(n4250), .I2(\useone/round_flag[5] ), 
            .I3(n1191_2), .O(n3527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6413.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6414 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[2] ), 
            .O(n4254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6414.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6415 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[4] ), 
            .I2(n4254), .I3(\useone/round_flag[0] ), .O(n4255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha73f */ ;
    defparam LUT__6415.LUTMASK = 16'ha73f;
    EFX_LUT4 LUT__6416 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[0] ), .O(n4256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8a7f */ ;
    defparam LUT__6416.LUTMASK = 16'h8a7f;
    EFX_LUT4 LUT__6417 (.I0(n4229), .I1(\useone/round_flag[1] ), .I2(n4256), 
            .O(n4257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__6417.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__6418 (.I0(n4257), .I1(n4255), .I2(\useone/round_flag[5] ), 
            .I3(n1191_2), .O(n3530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6418.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6419 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[5] ), .O(n4258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3c5 */ ;
    defparam LUT__6419.LUTMASK = 16'ha3c5;
    EFX_LUT4 LUT__6420 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[5] ), .O(n4259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1001 */ ;
    defparam LUT__6420.LUTMASK = 16'h1001;
    EFX_LUT4 LUT__6421 (.I0(\useone/round_flag[4] ), .I1(n4258), .I2(n4259), 
            .I3(\useone/round_flag[0] ), .O(n4260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6421.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6422 (.I0(n4228), .I1(\useone/round_flag[5] ), .I2(\useone/round_flag[4] ), 
            .I3(\useone/round_flag[2] ), .O(n4261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00b2 */ ;
    defparam LUT__6422.LUTMASK = 16'h00b2;
    EFX_LUT4 LUT__6423 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[5] ), .O(n4262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6100 */ ;
    defparam LUT__6423.LUTMASK = 16'h6100;
    EFX_LUT4 LUT__6424 (.I0(n4261), .I1(n4262), .I2(\useone/round_flag[0] ), 
            .I3(n4260), .O(n4263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f1 */ ;
    defparam LUT__6424.LUTMASK = 16'h00f1;
    EFX_LUT4 LUT__6425 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[5] ), 
            .O(n4264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6425.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6426 (.I0(\useone/round_flag[3] ), .I1(n4264), .I2(\useone/round_flag[0] ), 
            .I3(n4220), .O(n4265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0bb */ ;
    defparam LUT__6426.LUTMASK = 16'hb0bb;
    EFX_LUT4 LUT__6427 (.I0(n4265), .I1(n3943), .I2(n4263), .I3(n1191_2), 
            .O(n3533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6427.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6428 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[0] ), 
            .O(n4266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6428.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6429 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[4] ), 
            .I2(n3944), .I3(\useone/round_flag[1] ), .O(n4267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__6429.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__6430 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .I2(n4221), .I3(\useone/round_flag[4] ), .O(n4268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fab */ ;
    defparam LUT__6430.LUTMASK = 16'h0fab;
    EFX_LUT4 LUT__6431 (.I0(n3920), .I1(n4267), .I2(n4268), .I3(n4224), 
            .O(n4269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb000 */ ;
    defparam LUT__6431.LUTMASK = 16'hb000;
    EFX_LUT4 LUT__6432 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[0] ), .O(n4270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hba5d */ ;
    defparam LUT__6432.LUTMASK = 16'hba5d;
    EFX_LUT4 LUT__6433 (.I0(n4270), .I1(n3911), .I2(\useone/round_flag[4] ), 
            .I3(n4240), .O(n4271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6433.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6434 (.I0(n4220), .I1(n4266), .I2(n4269), .I3(n4271), 
            .O(n3536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__6434.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__6435 (.I0(\useone/round_flag[2] ), .I1(n3944), .I2(n4224), 
            .O(n4272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6435.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6436 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[4] ), .O(n4273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h384f */ ;
    defparam LUT__6436.LUTMASK = 16'h384f;
    EFX_LUT4 LUT__6437 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[2] ), .O(n4274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc07d */ ;
    defparam LUT__6437.LUTMASK = 16'hc07d;
    EFX_LUT4 LUT__6438 (.I0(n4274), .I1(n4273), .I2(\useone/round_flag[1] ), 
            .O(n4275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6438.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6439 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[0] ), .O(n4276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e03 */ ;
    defparam LUT__6439.LUTMASK = 16'h7e03;
    EFX_LUT4 LUT__6440 (.I0(n4276), .I1(n4227), .I2(n4275), .I3(n4272), 
            .O(n3539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f44 */ ;
    defparam LUT__6440.LUTMASK = 16'h4f44;
    EFX_LUT4 LUT__6441 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[4] ), .O(n4277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0017 */ ;
    defparam LUT__6441.LUTMASK = 16'h0017;
    EFX_LUT4 LUT__6442 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[1] ), .O(n4278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3ffd */ ;
    defparam LUT__6442.LUTMASK = 16'h3ffd;
    EFX_LUT4 LUT__6443 (.I0(n4237), .I1(n4278), .I2(\useone/round_flag[0] ), 
            .O(n4279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7c7c */ ;
    defparam LUT__6443.LUTMASK = 16'h7c7c;
    EFX_LUT4 LUT__6444 (.I0(\useone/round_flag[4] ), .I1(n4277), .I2(n4224), 
            .I3(n4279), .O(n4280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__6444.LUTMASK = 16'he000;
    EFX_LUT4 LUT__6445 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[2] ), 
            .O(n4281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6445.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6446 (.I0(\useone/round_flag[4] ), .I1(n3950), .I2(\useone/round_flag[0] ), 
            .I3(\useone/round_flag[2] ), .O(n4282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h87b8 */ ;
    defparam LUT__6446.LUTMASK = 16'h87b8;
    EFX_LUT4 LUT__6447 (.I0(n4281), .I1(n4282), .I2(\useone/round_flag[1] ), 
            .I3(n4240), .O(n4283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3500 */ ;
    defparam LUT__6447.LUTMASK = 16'h3500;
    EFX_LUT4 LUT__6448 (.I0(\useone/round_flag[4] ), .I1(n3944), .I2(n4283), 
            .I3(n4280), .O(n3542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0 */ ;
    defparam LUT__6448.LUTMASK = 16'hffe0;
    EFX_LUT4 LUT__6449 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[3] ), .O(n4284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e0d */ ;
    defparam LUT__6449.LUTMASK = 16'h3e0d;
    EFX_LUT4 LUT__6450 (.I0(n3931), .I1(n3910), .I2(n4284), .I3(\useone/round_flag[5] ), 
            .O(n4285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0bb */ ;
    defparam LUT__6450.LUTMASK = 16'hf0bb;
    EFX_LUT4 LUT__6451 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[5] ), .I3(\useone/round_flag[1] ), .O(n4286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h573c */ ;
    defparam LUT__6451.LUTMASK = 16'h573c;
    EFX_LUT4 LUT__6452 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .O(n4287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__6452.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__6453 (.I0(n3954), .I1(\useone/round_flag[5] ), .I2(n4287), 
            .I3(n4266), .O(n4288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6453.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6454 (.I0(\useone/round_flag[0] ), .I1(n4286), .I2(n4288), 
            .I3(n1191_2), .O(n4289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__6454.LUTMASK = 16'he000;
    EFX_LUT4 LUT__6455 (.I0(n4285), .I1(n1191_2), .I2(n4289), .I3(\useone/round_flag[4] ), 
            .O(n3545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf044 */ ;
    defparam LUT__6455.LUTMASK = 16'hf044;
    EFX_LUT4 LUT__6456 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8a3 */ ;
    defparam LUT__6456.LUTMASK = 16'hf8a3;
    EFX_LUT4 LUT__6457 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[2] ), 
            .I2(n4290), .O(n4291)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__6457.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__6458 (.I0(\useone/round_flag[0] ), .I1(n3910), .I2(\useone/round_flag[1] ), 
            .O(n4292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__6458.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__6459 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[2] ), 
            .O(n4293)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6459.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6460 (.I0(n4293), .I1(\useone/round_flag[0] ), .I2(n4287), 
            .I3(\useone/round_flag[5] ), .O(n4294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6460.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6461 (.I0(n4292), .I1(n3935), .I2(n4226), .I3(n4294), 
            .O(n4295)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6461.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6462 (.I0(n4291), .I1(\useone/round_flag[5] ), .I2(n4295), 
            .I3(n1191_2), .O(n3548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6462.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6463 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[4] ), .O(n4296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h70cf */ ;
    defparam LUT__6463.LUTMASK = 16'h70cf;
    EFX_LUT4 LUT__6464 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[3] ), .I3(n4296), .O(n4297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfd03 */ ;
    defparam LUT__6464.LUTMASK = 16'hfd03;
    EFX_LUT4 LUT__6465 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[0] ), 
            .O(n4298)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6465.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6466 (.I0(n4298), .I1(n3920), .I2(n3953), .O(n4299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6466.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6467 (.I0(n3932), .I1(n3937), .I2(\useone/round_flag[3] ), 
            .I3(n4299), .O(n4300)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6467.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6468 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .O(n4301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6468.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6469 (.I0(n4220), .I1(n4301), .I2(n4221), .I3(n4224), 
            .O(n4302)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6469.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6470 (.I0(n4300), .I1(n4240), .I2(n4297), .I3(n4302), 
            .O(n3551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__6470.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__6471 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[2] ), .O(n4303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8cf */ ;
    defparam LUT__6471.LUTMASK = 16'hf8cf;
    EFX_LUT4 LUT__6472 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4304)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6e8f */ ;
    defparam LUT__6472.LUTMASK = 16'h6e8f;
    EFX_LUT4 LUT__6473 (.I0(\useone/round_flag[3] ), .I1(n4304), .I2(n4224), 
            .O(n4305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__6473.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__6474 (.I0(n4254), .I1(n3944), .I2(n4248), .I3(\useone/round_flag[4] ), 
            .O(n4306)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6474.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6475 (.I0(\useone/round_flag[0] ), .I1(n3910), .I2(n4306), 
            .I3(n4240), .O(n4307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6475.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6476 (.I0(n4303), .I1(\useone/round_flag[0] ), .I2(n4305), 
            .I3(n4307), .O(n3554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffb0 */ ;
    defparam LUT__6476.LUTMASK = 16'hffb0;
    EFX_LUT4 LUT__6477 (.I0(n3925), .I1(n3937), .I2(n3909), .I3(\useone/round_flag[3] ), 
            .O(n4308)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heef0 */ ;
    defparam LUT__6477.LUTMASK = 16'heef0;
    EFX_LUT4 LUT__6478 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[0] ), .O(n4309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h83dc */ ;
    defparam LUT__6478.LUTMASK = 16'h83dc;
    EFX_LUT4 LUT__6479 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[0] ), .O(n4310)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hadc3 */ ;
    defparam LUT__6479.LUTMASK = 16'hadc3;
    EFX_LUT4 LUT__6480 (.I0(n4310), .I1(n4309), .I2(\useone/round_flag[5] ), 
            .I3(\useone/round_flag[4] ), .O(n4311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__6480.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__6481 (.I0(n4308), .I1(n4264), .I2(n4311), .I3(n1191_2), 
            .O(n3557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6481.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6482 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[1] ), .O(n4312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2cd7 */ ;
    defparam LUT__6482.LUTMASK = 16'h2cd7;
    EFX_LUT4 LUT__6483 (.I0(\useone/round_flag[4] ), .I1(n4312), .I2(n3906), 
            .O(n4313)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6483.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6484 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[3] ), .O(n4314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8a3f */ ;
    defparam LUT__6484.LUTMASK = 16'h8a3f;
    EFX_LUT4 LUT__6485 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[3] ), .O(n4315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb5f3 */ ;
    defparam LUT__6485.LUTMASK = 16'hb5f3;
    EFX_LUT4 LUT__6486 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[5] ), .O(n4316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6486.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6487 (.I0(n4315), .I1(n4314), .I2(\useone/round_flag[1] ), 
            .I3(n4316), .O(n4317)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha300 */ ;
    defparam LUT__6487.LUTMASK = 16'ha300;
    EFX_LUT4 LUT__6488 (.I0(\useone/round_flag[5] ), .I1(n4313), .I2(n4317), 
            .I3(n1191_2), .O(n3560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__6488.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__6489 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[1] ), .O(n4318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h45f3 */ ;
    defparam LUT__6489.LUTMASK = 16'h45f3;
    EFX_LUT4 LUT__6490 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[2] ), .O(n4319)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he1ae */ ;
    defparam LUT__6490.LUTMASK = 16'he1ae;
    EFX_LUT4 LUT__6491 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[0] ), .O(n4320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7c45 */ ;
    defparam LUT__6491.LUTMASK = 16'h7c45;
    EFX_LUT4 LUT__6492 (.I0(n4320), .I1(n4319), .I2(\useone/round_flag[4] ), 
            .I3(n4224), .O(n4321)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6492.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6493 (.I0(n4318), .I1(n4227), .I2(n4321), .O(n3563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__6493.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__6494 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[3] ), .O(n4322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcad8 */ ;
    defparam LUT__6494.LUTMASK = 16'hcad8;
    EFX_LUT4 LUT__6495 (.I0(\useone/round_flag[0] ), .I1(n3910), .I2(\useone/round_flag[4] ), 
            .I3(n4322), .O(n4323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f73 */ ;
    defparam LUT__6495.LUTMASK = 16'h0f73;
    EFX_LUT4 LUT__6496 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[2] ), .O(n4324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__6496.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__6497 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[0] ), 
            .I2(n4324), .I3(\useone/round_flag[4] ), .O(n4325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcdf0 */ ;
    defparam LUT__6497.LUTMASK = 16'hcdf0;
    EFX_LUT4 LUT__6498 (.I0(\useone/round_flag[3] ), .I1(n3902), .I2(n4325), 
            .I3(\useone/round_flag[5] ), .O(n4326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__6498.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__6499 (.I0(\useone/round_flag[5] ), .I1(n4323), .I2(n4326), 
            .I3(n1191_2), .O(n3566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__6499.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__6500 (.I0(\useone/round_flag[4] ), .I1(n4287), .I2(n4229), 
            .O(n4327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6500.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6501 (.I0(n3902), .I1(n4252), .I2(\useone/round_flag[0] ), 
            .I3(\useone/round_flag[3] ), .O(n4328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he00e */ ;
    defparam LUT__6501.LUTMASK = 16'he00e;
    EFX_LUT4 LUT__6502 (.I0(n4327), .I1(\useone/round_flag[0] ), .I2(n4328), 
            .I3(\useone/round_flag[5] ), .O(n4329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__6502.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__6503 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__6503.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__6504 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb200 */ ;
    defparam LUT__6504.LUTMASK = 16'hb200;
    EFX_LUT4 LUT__6505 (.I0(n4331), .I1(n4330), .I2(\useone/round_flag[2] ), 
            .I3(\useone/round_flag[3] ), .O(n4332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6505.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6506 (.I0(\useone/round_flag[3] ), .I1(n3943), .I2(n4226), 
            .I3(n4332), .O(n4333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__6506.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__6507 (.I0(n4333), .I1(n4329), .I2(n1191_2), .O(n3569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__6507.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__6508 (.I0(n4264), .I1(n1191_2), .O(n4334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6508.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6509 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[0] ), .O(n4335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbec0 */ ;
    defparam LUT__6509.LUTMASK = 16'hbec0;
    EFX_LUT4 LUT__6510 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[1] ), .O(n4336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf03b */ ;
    defparam LUT__6510.LUTMASK = 16'hf03b;
    EFX_LUT4 LUT__6511 (.I0(n4336), .I1(n3911), .I2(\useone/round_flag[4] ), 
            .I3(n4240), .O(n4337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5c00 */ ;
    defparam LUT__6511.LUTMASK = 16'h5c00;
    EFX_LUT4 LUT__6512 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[3] ), .O(n4338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4dbe */ ;
    defparam LUT__6512.LUTMASK = 16'h4dbe;
    EFX_LUT4 LUT__6513 (.I0(n4338), .I1(n1191_2), .I2(\useone/round_flag[4] ), 
            .I3(\useone/round_flag[5] ), .O(n4339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6513.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6514 (.I0(n4335), .I1(n4334), .I2(n4337), .I3(n4339), 
            .O(n3572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff8 */ ;
    defparam LUT__6514.LUTMASK = 16'hfff8;
    EFX_LUT4 LUT__6515 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[4] ), .O(n4340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3fe */ ;
    defparam LUT__6515.LUTMASK = 16'hd3fe;
    EFX_LUT4 LUT__6516 (.I0(n4241), .I1(\useone/round_flag[2] ), .I2(\useone/round_flag[4] ), 
            .O(n4341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6516.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6517 (.I0(\useone/round_flag[1] ), .I1(n4340), .I2(n4341), 
            .O(n4342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__6517.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6518 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[3] ), .O(n4343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9d78 */ ;
    defparam LUT__6518.LUTMASK = 16'h9d78;
    EFX_LUT4 LUT__6519 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[0] ), .O(n4344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6519.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6520 (.I0(n4248), .I1(n4220), .I2(n4221), .I3(n4344), 
            .O(n4345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6520.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6521 (.I0(\useone/round_flag[2] ), .I1(n4343), .I2(n4224), 
            .I3(n4345), .O(n4346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__6521.LUTMASK = 16'he000;
    EFX_LUT4 LUT__6522 (.I0(n4342), .I1(n4240), .I2(n4346), .O(n3575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__6522.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__6523 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[2] ), .O(n4347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha8d3 */ ;
    defparam LUT__6523.LUTMASK = 16'ha8d3;
    EFX_LUT4 LUT__6524 (.I0(n3910), .I1(\useone/round_flag[4] ), .I2(n4347), 
            .O(n4348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd3d3 */ ;
    defparam LUT__6524.LUTMASK = 16'hd3d3;
    EFX_LUT4 LUT__6525 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[3] ), .O(n4349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h533d */ ;
    defparam LUT__6525.LUTMASK = 16'h533d;
    EFX_LUT4 LUT__6526 (.I0(n4224), .I1(n4349), .I2(\useone/round_flag[4] ), 
            .O(n4350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6526.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6527 (.I0(\useone/round_flag[0] ), .I1(n4287), .I2(n4281), 
            .I3(n4334), .O(n4351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6527.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6528 (.I0(n4348), .I1(n4240), .I2(n4350), .I3(n4351), 
            .O(n3578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__6528.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__6529 (.I0(n4224), .I1(\useone/round_flag[4] ), .O(n4352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6529.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6530 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[2] ), .O(n4353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h73e5 */ ;
    defparam LUT__6530.LUTMASK = 16'h73e5;
    EFX_LUT4 LUT__6531 (.I0(n4228), .I1(n3954), .I2(\useone/round_flag[0] ), 
            .I3(n4334), .O(n4354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e00 */ ;
    defparam LUT__6531.LUTMASK = 16'h3e00;
    EFX_LUT4 LUT__6532 (.I0(\useone/round_flag[2] ), .I1(\useone/n46233 ), 
            .I2(n4248), .I3(\useone/round_flag[4] ), .O(n4355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__6532.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__6533 (.I0(\useone/round_flag[4] ), .I1(n3911), .I2(n4355), 
            .I3(n4240), .O(n4356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__6533.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__6534 (.I0(n4353), .I1(n4352), .I2(n4354), .I3(n4356), 
            .O(n3581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfff4 */ ;
    defparam LUT__6534.LUTMASK = 16'hfff4;
    EFX_LUT4 LUT__6535 (.I0(\useone/round_flag[4] ), .I1(n3911), .O(n4357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6535.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6536 (.I0(n3955), .I1(n4301), .I2(n4236), .I3(\useone/round_flag[4] ), 
            .O(n4358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6536.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6537 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[4] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[1] ), .O(n4359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ecf */ ;
    defparam LUT__6537.LUTMASK = 16'h5ecf;
    EFX_LUT4 LUT__6538 (.I0(n4281), .I1(\useone/round_flag[4] ), .I2(\useone/round_flag[0] ), 
            .I3(\useone/round_flag[1] ), .O(n4360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h57c5 */ ;
    defparam LUT__6538.LUTMASK = 16'h57c5;
    EFX_LUT4 LUT__6539 (.I0(\useone/round_flag[2] ), .I1(n4359), .I2(n4360), 
            .I3(n4224), .O(n4361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__6539.LUTMASK = 16'he000;
    EFX_LUT4 LUT__6540 (.I0(n4358), .I1(n4357), .I2(n4240), .I3(n4361), 
            .O(n3584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hffe0 */ ;
    defparam LUT__6540.LUTMASK = 16'hffe0;
    EFX_LUT4 LUT__6541 (.I0(n4344), .I1(n3944), .I2(\useone/round_flag[2] ), 
            .O(n4362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6541.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6542 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[4] ), .O(n4363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__6542.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__6543 (.I0(n4254), .I1(n3920), .I2(n4363), .I3(\useone/round_flag[5] ), 
            .O(n4364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6543.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6544 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[1] ), .O(n4365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3edf */ ;
    defparam LUT__6544.LUTMASK = 16'h3edf;
    EFX_LUT4 LUT__6545 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[3] ), .O(n4366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6545.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6546 (.I0(n4254), .I1(\useone/round_flag[4] ), .I2(n4366), 
            .I3(\useone/round_flag[5] ), .O(n4367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__6546.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__6547 (.I0(\useone/round_flag[2] ), .I1(n4365), .I2(n4367), 
            .O(n4368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6547.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6548 (.I0(n4364), .I1(n4362), .I2(n4368), .I3(n1191_2), 
            .O(n3587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6548.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6549 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[1] ), .O(n4369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h30d7 */ ;
    defparam LUT__6549.LUTMASK = 16'h30d7;
    EFX_LUT4 LUT__6550 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[0] ), .I3(n4281), .O(n4370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc8bf */ ;
    defparam LUT__6550.LUTMASK = 16'hc8bf;
    EFX_LUT4 LUT__6551 (.I0(n3937), .I1(\useone/round_flag[0] ), .I2(\useone/round_flag[5] ), 
            .I3(\useone/round_flag[3] ), .O(n4371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b00 */ ;
    defparam LUT__6551.LUTMASK = 16'h2b00;
    EFX_LUT4 LUT__6552 (.I0(n4371), .I1(\useone/round_flag[4] ), .I2(n4370), 
            .O(n4372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6552.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6553 (.I0(\useone/round_flag[3] ), .I1(n4254), .I2(\useone/round_flag[4] ), 
            .I3(n1191_2), .O(n4373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6553.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6554 (.I0(n3955), .I1(\useone/round_flag[5] ), .I2(n1191_2), 
            .I3(n4373), .O(n4374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__6554.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__6555 (.I0(n4369), .I1(n4264), .I2(n4372), .I3(n4374), 
            .O(n3590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000b */ ;
    defparam LUT__6555.LUTMASK = 16'h000b;
    EFX_LUT4 LUT__6556 (.I0(n4228), .I1(n3932), .I2(\useone/round_flag[5] ), 
            .O(n4375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6556.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6557 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .I3(n3950), .O(n4376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd5dc */ ;
    defparam LUT__6557.LUTMASK = 16'hd5dc;
    EFX_LUT4 LUT__6558 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[0] ), .O(n4377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h730f */ ;
    defparam LUT__6558.LUTMASK = 16'h730f;
    EFX_LUT4 LUT__6559 (.I0(\useone/round_flag[4] ), .I1(n4248), .I2(n4266), 
            .O(n4378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4141 */ ;
    defparam LUT__6559.LUTMASK = 16'h4141;
    EFX_LUT4 LUT__6560 (.I0(\useone/round_flag[4] ), .I1(n4377), .I2(n4378), 
            .I3(n4224), .O(n4379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6560.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6561 (.I0(n4376), .I1(n4373), .I2(n4375), .I3(n4379), 
            .O(n3593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff80 */ ;
    defparam LUT__6561.LUTMASK = 16'hff80;
    EFX_LUT4 LUT__6562 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[2] ), .O(n4380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6562.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6563 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[0] ), .O(n4381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he800 */ ;
    defparam LUT__6563.LUTMASK = 16'he800;
    EFX_LUT4 LUT__6564 (.I0(\useone/round_flag[3] ), .I1(n4293), .I2(\useone/round_flag[5] ), 
            .O(n4382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6564.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6565 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heb00 */ ;
    defparam LUT__6565.LUTMASK = 16'heb00;
    EFX_LUT4 LUT__6566 (.I0(n3931), .I1(n4383), .O(n4384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6566.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6567 (.I0(\useone/round_flag[5] ), .I1(n4384), .I2(n3955), 
            .I3(n1191_2), .O(n4385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6567.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6568 (.I0(n4381), .I1(n4380), .I2(n4382), .I3(n4385), 
            .O(n3596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6568.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6569 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[3] ), .O(n4386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf8a3 */ ;
    defparam LUT__6569.LUTMASK = 16'hf8a3;
    EFX_LUT4 LUT__6570 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7ffc */ ;
    defparam LUT__6570.LUTMASK = 16'h7ffc;
    EFX_LUT4 LUT__6571 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[0] ), .I3(\useone/round_flag[1] ), .O(n4388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h83fa */ ;
    defparam LUT__6571.LUTMASK = 16'h83fa;
    EFX_LUT4 LUT__6572 (.I0(n4387), .I1(\useone/round_flag[3] ), .I2(n4388), 
            .I3(\useone/round_flag[5] ), .O(n4389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6572.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6573 (.I0(n4386), .I1(n4226), .I2(n4374), .I3(n4389), 
            .O(n3599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6573.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6574 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[2] ), .O(n4390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc3fd */ ;
    defparam LUT__6574.LUTMASK = 16'hc3fd;
    EFX_LUT4 LUT__6575 (.I0(n3909), .I1(\useone/round_flag[3] ), .I2(n4390), 
            .I3(\useone/round_flag[4] ), .O(n4391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h70cc */ ;
    defparam LUT__6575.LUTMASK = 16'h70cc;
    EFX_LUT4 LUT__6576 (.I0(\useone/round_flag[0] ), .I1(n4391), .I2(\useone/round_flag[4] ), 
            .I3(n3943), .O(n4392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0dc3 */ ;
    defparam LUT__6576.LUTMASK = 16'h0dc3;
    EFX_LUT4 LUT__6577 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[3] ), .O(n4393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4b00 */ ;
    defparam LUT__6577.LUTMASK = 16'h4b00;
    EFX_LUT4 LUT__6578 (.I0(n3925), .I1(n3902), .I2(n4220), .O(n4394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6578.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6579 (.I0(n4394), .I1(n4393), .I2(n4373), .I3(n4224), 
            .O(n4395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6579.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6580 (.I0(\useone/round_flag[5] ), .I1(n4392), .I2(n4395), 
            .O(n3602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6580.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6581 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[1] ), .O(n4396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd274 */ ;
    defparam LUT__6581.LUTMASK = 16'hd274;
    EFX_LUT4 LUT__6582 (.I0(n4396), .I1(n3911), .I2(\useone/round_flag[4] ), 
            .O(n4397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'ha3a3 */ ;
    defparam LUT__6582.LUTMASK = 16'ha3a3;
    EFX_LUT4 LUT__6583 (.I0(n4254), .I1(\useone/round_flag[0] ), .I2(\useone/round_flag[3] ), 
            .I3(\useone/round_flag[4] ), .O(n4398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hafdc */ ;
    defparam LUT__6583.LUTMASK = 16'hafdc;
    EFX_LUT4 LUT__6584 (.I0(n3937), .I1(\useone/round_flag[3] ), .I2(\useone/round_flag[0] ), 
            .I3(n4398), .O(n4399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__6584.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__6585 (.I0(n4399), .I1(n4397), .I2(\useone/round_flag[5] ), 
            .I3(n1191_2), .O(n3605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5300 */ ;
    defparam LUT__6585.LUTMASK = 16'h5300;
    EFX_LUT4 LUT__6586 (.I0(\useone/round_flag[1] ), .I1(n3918), .O(n4400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6586.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6587 (.I0(n3933), .I1(n3923), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[2] ), .O(n4401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5333 */ ;
    defparam LUT__6587.LUTMASK = 16'h5333;
    EFX_LUT4 LUT__6588 (.I0(\useone/round_flag[5] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[3] ), .O(n4402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6588.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6589 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[4] ), .O(n4403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3001 */ ;
    defparam LUT__6589.LUTMASK = 16'h3001;
    EFX_LUT4 LUT__6590 (.I0(n3927), .I1(\useone/round_flag[1] ), .I2(n3917), 
            .I3(\useone/round_flag[2] ), .O(n4404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6590.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6591 (.I0(n4403), .I1(n4402), .I2(n4404), .I3(n3938), 
            .O(n4405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6591.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6592 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .O(n4406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6592.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6593 (.I0(n3901), .I1(n4406), .O(n4407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6593.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6594 (.I0(n3917), .I1(n3937), .O(n4408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6594.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6595 (.I0(n3924), .I1(n4254), .I2(n4407), .I3(n4408), 
            .O(n4409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6595.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6596 (.I0(n4400), .I1(n4401), .I2(n4405), .I3(n4409), 
            .O(n3608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6596.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6597 (.I0(n3927), .I1(n3918), .I2(\useone/round_flag[2] ), 
            .O(n4410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6597.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6598 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[4] ), 
            .O(n4411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6598.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6599 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[5] ), .O(n4412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6599.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6600 (.I0(n4411), .I1(n4412), .I2(n3943), .O(n4413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6600.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6601 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[1] ), .O(n4414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6601.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6602 (.I0(n4414), .I1(n3924), .I2(\useone/round_flag[2] ), 
            .I3(\useone/round_flag[0] ), .O(n4415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6602.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6603 (.I0(\useone/round_flag[1] ), .I1(n4410), .I2(n4413), 
            .I3(n4415), .O(n4416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000e */ ;
    defparam LUT__6603.LUTMASK = 16'h000e;
    EFX_LUT4 LUT__6604 (.I0(n3913), .I1(n3901), .I2(n3917), .I3(n3953), 
            .O(n4417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6604.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6605 (.I0(n3912), .I1(n3955), .I2(n3904), .I3(n4417), 
            .O(n4418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6605.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6606 (.I0(\useone/round_flag[0] ), .I1(n3902), .I2(n3923), 
            .O(n4419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6606.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6607 (.I0(n3935), .I1(n3927), .O(n4420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6607.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6608 (.I0(n3905), .I1(n3924), .I2(\useone/round_flag[2] ), 
            .I3(\useone/round_flag[1] ), .O(n4421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6608.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6609 (.I0(n4419), .I1(n4420), .I2(n4421), .O(n4422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__6609.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__6610 (.I0(n3923), .I1(n3917), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[2] ), .O(n4423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0a0c */ ;
    defparam LUT__6610.LUTMASK = 16'h0a0c;
    EFX_LUT4 LUT__6611 (.I0(n3912), .I1(n3949), .I2(n3924), .I3(n3902), 
            .O(n4424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6611.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6612 (.I0(n4423), .I1(n4424), .O(n4425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6612.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6613 (.I0(n4416), .I1(n4418), .I2(n4422), .I3(n4425), 
            .O(n3611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6613.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6614 (.I0(n3903), .I1(n3917), .I2(\useone/n46233 ), 
            .I3(\useone/round_flag[2] ), .O(n4426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6614.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6615 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(n3901), .O(n4427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1400 */ ;
    defparam LUT__6615.LUTMASK = 16'h1400;
    EFX_LUT4 LUT__6616 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .I3(n3927), .O(n4428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9e00 */ ;
    defparam LUT__6616.LUTMASK = 16'h9e00;
    EFX_LUT4 LUT__6617 (.I0(n3903), .I1(n4266), .I2(n3937), .I3(n3918), 
            .O(n4429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f */ ;
    defparam LUT__6617.LUTMASK = 16'h035f;
    EFX_LUT4 LUT__6618 (.I0(n3933), .I1(n3917), .I2(n4254), .O(n4430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6618.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6619 (.I0(n4419), .I1(n4428), .I2(n4430), .I3(n4429), 
            .O(n4431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6619.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6620 (.I0(n3923), .I1(n3933), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[2] ), .O(n4432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6620.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6621 (.I0(n3935), .I1(n3928), .I2(n3924), .I3(n4432), 
            .O(n4433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6621.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6622 (.I0(n4426), .I1(n4427), .I2(n4431), .I3(n4433), 
            .O(n3614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefff */ ;
    defparam LUT__6622.LUTMASK = 16'hefff;
    EFX_LUT4 LUT__6623 (.I0(n4254), .I1(n3917), .I2(n3901), .I3(n4221), 
            .O(n4434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f */ ;
    defparam LUT__6623.LUTMASK = 16'h035f;
    EFX_LUT4 LUT__6624 (.I0(n3934), .I1(n4420), .I2(n4434), .O(n4435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6624.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6625 (.I0(\useone/round_flag[0] ), .I1(n3918), .I2(n3903), 
            .I3(n4254), .O(n4436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6625.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6626 (.I0(n3927), .I1(n4221), .I2(n3923), .I3(n3902), 
            .O(n4437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6626.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6627 (.I0(n3912), .I1(n4242), .I2(n3918), .I3(n3937), 
            .O(n4438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6627.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6628 (.I0(n4436), .I1(n4437), .I2(n4438), .O(n4439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6628.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6629 (.I0(n3924), .I1(n3902), .O(n4440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6629.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6630 (.I0(n3900), .I1(n3903), .I2(n3918), .I3(n3932), 
            .O(n4441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6630.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6631 (.I0(n4440), .I1(n4423), .I2(n4441), .O(n4442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6631.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6632 (.I0(n3916), .I1(n4435), .I2(n4439), .I3(n4442), 
            .O(n3617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6632.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6633 (.I0(n3901), .I1(\useone/round_flag[0] ), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[2] ), .O(n4443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he00e */ ;
    defparam LUT__6633.LUTMASK = 16'he00e;
    EFX_LUT4 LUT__6634 (.I0(n3924), .I1(n3923), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[0] ), .O(n4444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf100 */ ;
    defparam LUT__6634.LUTMASK = 16'hf100;
    EFX_LUT4 LUT__6635 (.I0(n4254), .I1(n3924), .I2(n4443), .I3(n4444), 
            .O(n4445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f4 */ ;
    defparam LUT__6635.LUTMASK = 16'h00f4;
    EFX_LUT4 LUT__6636 (.I0(\useone/round_flag[6] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[4] ), .O(n4446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6636.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6637 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[3] ), 
            .I2(n4446), .I3(n3931), .O(n4447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000 */ ;
    defparam LUT__6637.LUTMASK = 16'h6000;
    EFX_LUT4 LUT__6638 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[5] ), .O(n4448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b2b */ ;
    defparam LUT__6638.LUTMASK = 16'h2b2b;
    EFX_LUT4 LUT__6639 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[3] ), .O(n4449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6639.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6640 (.I0(n4448), .I1(n4449), .I2(n4254), .I3(n3903), 
            .O(n4450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6640.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6641 (.I0(\useone/round_flag[2] ), .I1(n3903), .I2(n4447), 
            .I3(n4450), .O(n4451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6641.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6642 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[1] ), .O(n4452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__6642.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__6643 (.I0(n3933), .I1(n4452), .I2(n3914), .I3(n3927), 
            .O(n4453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6643.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6644 (.I0(n4445), .I1(n3929), .I2(n4451), .I3(n4453), 
            .O(n3620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefff */ ;
    defparam LUT__6644.LUTMASK = 16'hefff;
    EFX_LUT4 LUT__6645 (.I0(n3925), .I1(n3917), .I2(n3924), .O(n4454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6645.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6646 (.I0(n3923), .I1(\useone/round_flag[0] ), .I2(n3901), 
            .I3(n3937), .O(n4455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6646.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6647 (.I0(\useone/round_flag[2] ), .I1(n4454), .I2(n4455), 
            .O(n4456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__6647.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6648 (.I0(n4242), .I1(n3912), .I2(n4408), .I3(n3936), 
            .O(n4457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6648.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6649 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[0] ), 
            .I2(n3910), .I3(\useone/round_flag[1] ), .O(n4458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbaf0 */ ;
    defparam LUT__6649.LUTMASK = 16'hbaf0;
    EFX_LUT4 LUT__6650 (.I0(\useone/round_flag[6] ), .I1(\useone/round_flag[5] ), 
            .O(n4459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6650.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6651 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[5] ), .O(n4460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbc00 */ ;
    defparam LUT__6651.LUTMASK = 16'hbc00;
    EFX_LUT4 LUT__6652 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[6] ), .O(n4461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__6652.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__6653 (.I0(n3954), .I1(\useone/round_flag[4] ), .I2(n4460), 
            .I3(n4461), .O(n4462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__6653.LUTMASK = 16'he000;
    EFX_LUT4 LUT__6654 (.I0(n4220), .I1(n4459), .I2(n4458), .I3(n4462), 
            .O(n4463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__6654.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__6655 (.I0(n3909), .I1(n3924), .I2(n3918), .I3(\useone/round_flag[2] ), 
            .O(n4464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6655.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6656 (.I0(n4413), .I1(n4464), .O(n4465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6656.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6657 (.I0(n4456), .I1(n4457), .I2(n4463), .I3(n4465), 
            .O(n3623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6657.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6658 (.I0(n3924), .I1(\useone/round_flag[0] ), .I2(n3917), 
            .I3(n3902), .O(n4466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__6658.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__6659 (.I0(n3927), .I1(n3902), .I2(n3935), .I3(n3923), 
            .O(n4467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6659.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6660 (.I0(n3923), .I1(n3949), .I2(n3909), .I3(n3924), 
            .O(n4468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6660.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6661 (.I0(n3923), .I1(n3937), .I2(n4467), .I3(n4468), 
            .O(n4469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__6661.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__6662 (.I0(\useone/round_flag[2] ), .I1(n4301), .I2(n3905), 
            .O(n4470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6662.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6663 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[4] ), 
            .I2(n4266), .I3(n4402), .O(n4471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9000 */ ;
    defparam LUT__6663.LUTMASK = 16'h9000;
    EFX_LUT4 LUT__6664 (.I0(n3924), .I1(n4452), .O(n4472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6664.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6665 (.I0(n3934), .I1(n4470), .I2(n4471), .I3(n4472), 
            .O(n4473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6665.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6666 (.I0(n3903), .I1(\useone/n46233 ), .I2(n4402), 
            .I3(n4221), .O(n4474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6666.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6667 (.I0(n3906), .I1(n3912), .I2(n4474), .O(n4475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__6667.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__6668 (.I0(n4466), .I1(n4469), .I2(n4473), .I3(n4475), 
            .O(n3626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6668.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6669 (.I0(n3923), .I1(\useone/round_flag[0] ), .I2(n3924), 
            .I3(\useone/round_flag[1] ), .O(n4476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__6669.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__6670 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[6] ), .I3(n3937), .O(n4477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6670.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6671 (.I0(n4266), .I1(n4477), .I2(n4476), .I3(n3927), 
            .O(n4478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heee0 */ ;
    defparam LUT__6671.LUTMASK = 16'heee0;
    EFX_LUT4 LUT__6672 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .O(n4479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6672.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6673 (.I0(n3923), .I1(n3913), .I2(n4479), .I3(n3933), 
            .O(n4480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6673.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6674 (.I0(n4400), .I1(n3927), .I2(n3932), .I3(n4480), 
            .O(n4481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__6674.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__6675 (.I0(n3901), .I1(n3914), .I2(n4446), .I3(n4242), 
            .O(n4482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6675.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6676 (.I0(n4221), .I1(n4412), .I2(n3902), .I3(n3901), 
            .O(n4483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6676.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6677 (.I0(n3927), .I1(n3943), .I2(n4482), .I3(n4483), 
            .O(n4484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__6677.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__6678 (.I0(n3918), .I1(n3914), .O(n4485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6678.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6679 (.I0(n4446), .I1(n3906), .O(n4486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6679.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6680 (.I0(n3913), .I1(n3924), .I2(n4485), .I3(n4486), 
            .O(n4487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6680.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6681 (.I0(n4478), .I1(n4481), .I2(n4484), .I3(n4487), 
            .O(n3629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6681.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6682 (.I0(n3927), .I1(n3901), .I2(\useone/round_flag[2] ), 
            .I3(n3909), .O(n4488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6682.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6683 (.I0(n4221), .I1(n3917), .I2(n4486), .I3(n4488), 
            .O(n4489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6683.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6684 (.I0(n3935), .I1(n3903), .O(n4490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6684.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6685 (.I0(n3949), .I1(n3923), .I2(n4490), .I3(n4440), 
            .O(n4491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6685.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6686 (.I0(\useone/round_flag[1] ), .I1(n3924), .I2(n3901), 
            .I3(\useone/round_flag[2] ), .O(n4492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__6686.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__6687 (.I0(n3907), .I1(n4408), .I2(n4420), .I3(n4492), 
            .O(n4493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6687.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6688 (.I0(n3914), .I1(n3903), .O(n4494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6688.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6689 (.I0(n3900), .I1(n4412), .O(n4495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6689.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6690 (.I0(\useone/round_flag[0] ), .I1(n3924), .I2(n3918), 
            .I3(n3952), .O(n4496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0bbb */ ;
    defparam LUT__6690.LUTMASK = 16'h0bbb;
    EFX_LUT4 LUT__6691 (.I0(n4423), .I1(n4494), .I2(n4495), .I3(n4496), 
            .O(n4497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6691.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6692 (.I0(n4489), .I1(n4491), .I2(n4493), .I3(n4497), 
            .O(n3632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6692.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6693 (.I0(n3923), .I1(n3937), .I2(n4466), .O(n4498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6693.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6694 (.I0(n3923), .I1(n3953), .I2(n3943), .I3(n3924), 
            .O(n4499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6694.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6695 (.I0(n3945), .I1(n3924), .I2(n3933), .I3(n4406), 
            .O(n4500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6695.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6696 (.I0(n4446), .I1(n4242), .I2(n3918), .I3(n4221), 
            .O(n4501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6696.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6697 (.I0(n4499), .I1(n4500), .I2(n4501), .O(n4502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6697.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6698 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .O(n4503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__6698.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__6699 (.I0(n3901), .I1(n4503), .O(n4504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6699.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6700 (.I0(n3927), .I1(n3943), .I2(n4490), .I3(n4504), 
            .O(n4505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6700.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6701 (.I0(n4457), .I1(n4498), .I2(n4502), .I3(n4505), 
            .O(n3635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6701.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6702 (.I0(\useone/round_flag[2] ), .I1(n3917), .I2(n3903), 
            .I3(\useone/round_flag[1] ), .O(n4506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__6702.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__6703 (.I0(n4506), .I1(\useone/round_flag[0] ), .O(n4507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6703.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6704 (.I0(n3923), .I1(n3914), .I2(n3917), .I3(n3913), 
            .O(n4508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6704.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6705 (.I0(n3903), .I1(n4468), .I2(n4254), .I3(n4508), 
            .O(n4509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f00 */ ;
    defparam LUT__6705.LUTMASK = 16'h4f00;
    EFX_LUT4 LUT__6706 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .O(n4510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6706.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6707 (.I0(\useone/round_flag[1] ), .I1(n3923), .I2(n3933), 
            .I3(n4510), .O(n4511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6707.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6708 (.I0(n3927), .I1(n3918), .I2(\useone/round_flag[2] ), 
            .I3(\useone/round_flag[0] ), .O(n4512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6708.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6709 (.I0(n3932), .I1(n3927), .I2(n3918), .I3(\useone/round_flag[1] ), 
            .O(n4513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__6709.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__6710 (.I0(n4511), .I1(n4512), .I2(n4513), .I3(n4499), 
            .O(n4514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6710.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6711 (.I0(n3924), .I1(n3917), .I2(n3902), .O(n4515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6711.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6712 (.I0(n3927), .I1(n3900), .O(n4516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6712.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6713 (.I0(n3934), .I1(n4427), .I2(n4515), .I3(n4516), 
            .O(n4517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6713.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6714 (.I0(n4507), .I1(n4509), .I2(n4514), .I3(n4517), 
            .O(n3638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6714.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6715 (.I0(n3927), .I1(n3903), .I2(\useone/round_flag[2] ), 
            .I3(n3923), .O(n4518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__6715.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__6716 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(n4412), .I3(n4518), .O(n4519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f8a */ ;
    defparam LUT__6716.LUTMASK = 16'h7f8a;
    EFX_LUT4 LUT__6717 (.I0(n3927), .I1(n4254), .I2(n4266), .I3(n3918), 
            .O(n4520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f */ ;
    defparam LUT__6717.LUTMASK = 16'h035f;
    EFX_LUT4 LUT__6718 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[3] ), .O(n4521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe3f */ ;
    defparam LUT__6718.LUTMASK = 16'hfe3f;
    EFX_LUT4 LUT__6719 (.I0(n3925), .I1(n4521), .I2(\useone/round_flag[5] ), 
            .I3(\useone/round_flag[6] ), .O(n4522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6719.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6720 (.I0(n4411), .I1(n4412), .I2(n4254), .O(n4523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6720.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6721 (.I0(n4404), .I1(n4523), .I2(n4492), .O(n4524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6721.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6722 (.I0(n4522), .I1(n4520), .I2(n4519), .I3(n4524), 
            .O(n3641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6722.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6723 (.I0(n3943), .I1(n3933), .I2(n3917), .I3(n3925), 
            .O(n4525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6723.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6724 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[0] ), 
            .I2(\useone/round_flag[2] ), .O(n4526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6724.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6725 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[2] ), .O(n4527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__6725.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6726 (.I0(n3905), .I1(n4527), .I2(n4526), .I3(n3901), 
            .O(n4528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__6726.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__6727 (.I0(\useone/n46233 ), .I1(n3918), .I2(n3903), 
            .I3(\useone/round_flag[2] ), .O(n4529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0fbb */ ;
    defparam LUT__6727.LUTMASK = 16'h0fbb;
    EFX_LUT4 LUT__6728 (.I0(n4525), .I1(n4528), .I2(n4529), .O(n4530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__6728.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__6729 (.I0(n4242), .I1(n4446), .I2(n4467), .O(n4531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__6729.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__6730 (.I0(n3917), .I1(n3928), .I2(n3918), .I3(n3902), 
            .O(n4532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6730.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6731 (.I0(n3912), .I1(n3906), .I2(n3923), .I3(n3902), 
            .O(n4533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6731.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6732 (.I0(n4532), .I1(n4533), .O(n4534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6732.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6733 (.I0(n4433), .I1(n4530), .I2(n4531), .I3(n4534), 
            .O(n3644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6733.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6734 (.I0(n3927), .I1(n3903), .I2(n3918), .I3(n3909), 
            .O(n4535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__6734.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__6735 (.I0(n3931), .I1(n3901), .I2(n4535), .I3(\useone/round_flag[2] ), 
            .O(n4536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6735.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6736 (.I0(n4254), .I1(n3927), .I2(n4266), .I3(n3917), 
            .O(n4537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0 */ ;
    defparam LUT__6736.LUTMASK = 16'hfac0;
    EFX_LUT4 LUT__6737 (.I0(n4400), .I1(n3933), .I2(n4510), .I3(n4537), 
            .O(n4538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__6737.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__6738 (.I0(n3949), .I1(n3924), .I2(n3901), .I3(n3914), 
            .O(n4539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h035f */ ;
    defparam LUT__6738.LUTMASK = 16'h035f;
    EFX_LUT4 LUT__6739 (.I0(n4419), .I1(n4539), .I2(n4468), .O(n4540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6739.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6740 (.I0(n4536), .I1(n4509), .I2(n4538), .I3(n4540), 
            .O(n3647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6740.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6741 (.I0(n3923), .I1(n3925), .I2(n3918), .I3(n3900), 
            .O(n4541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6741.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6742 (.I0(n3923), .I1(n3924), .I2(n4254), .I3(n4541), 
            .O(n4542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__6742.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__6743 (.I0(\useone/round_flag[5] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[3] ), .O(n4543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6743.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6744 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[4] ), .I3(n4543), .O(n4544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h2b00 */ ;
    defparam LUT__6744.LUTMASK = 16'h2b00;
    EFX_LUT4 LUT__6745 (.I0(n3933), .I1(n3902), .I2(n3918), .I3(n4510), 
            .O(n4545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6745.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6746 (.I0(n4447), .I1(n4544), .I2(n4545), .I3(n4437), 
            .O(n4546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6746.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6747 (.I0(n3923), .I1(n3945), .I2(n4254), .I3(n3901), 
            .O(n4547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6747.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6748 (.I0(n4523), .I1(n4525), .I2(n4547), .O(n4548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6748.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6749 (.I0(n4254), .I1(n3927), .I2(n3933), .I3(n3932), 
            .O(n4549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6749.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6750 (.I0(n4542), .I1(n4546), .I2(n4548), .I3(n4549), 
            .O(n3650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6750.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6751 (.I0(n4523), .I1(n4547), .O(n4550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6751.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6752 (.I0(n3927), .I1(n3923), .I2(\useone/round_flag[0] ), 
            .I3(\useone/round_flag[2] ), .O(n4551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1ff3 */ ;
    defparam LUT__6752.LUTMASK = 16'h1ff3;
    EFX_LUT4 LUT__6753 (.I0(\useone/round_flag[1] ), .I1(n4551), .I2(n4516), 
            .O(n4552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__6753.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__6754 (.I0(\useone/round_flag[4] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[0] ), .O(n4553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h15cf */ ;
    defparam LUT__6754.LUTMASK = 16'h15cf;
    EFX_LUT4 LUT__6755 (.I0(n4553), .I1(n4402), .I2(n4537), .O(n4554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6755.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6756 (.I0(n3917), .I1(\useone/round_flag[0] ), .I2(n3924), 
            .I3(n3902), .O(n4555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h15cf */ ;
    defparam LUT__6756.LUTMASK = 16'h15cf;
    EFX_LUT4 LUT__6757 (.I0(n4550), .I1(n4552), .I2(n4554), .I3(n4555), 
            .O(n3653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6757.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6758 (.I0(n3932), .I1(n4532), .I2(n4402), .I3(n4522), 
            .O(n4556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h007f */ ;
    defparam LUT__6758.LUTMASK = 16'h007f;
    EFX_LUT4 LUT__6759 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[3] ), .I3(\useone/round_flag[4] ), .O(n4557)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe8f */ ;
    defparam LUT__6759.LUTMASK = 16'hfe8f;
    EFX_LUT4 LUT__6760 (.I0(n4557), .I1(\useone/round_flag[0] ), .I2(n4459), 
            .I3(n4494), .O(n4558)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00ef */ ;
    defparam LUT__6760.LUTMASK = 16'h00ef;
    EFX_LUT4 LUT__6761 (.I0(\useone/round_flag[6] ), .I1(\useone/round_flag[3] ), 
            .O(n4559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6761.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6762 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[5] ), 
            .I2(\useone/round_flag[4] ), .I3(n4559), .O(n4560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6100 */ ;
    defparam LUT__6762.LUTMASK = 16'h6100;
    EFX_LUT4 LUT__6763 (.I0(\useone/round_flag[3] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[1] ), .O(n4561)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6763.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6764 (.I0(n4561), .I1(n3927), .I2(n3917), .I3(n4221), 
            .O(n4562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__6764.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__6765 (.I0(n4254), .I1(n4560), .I2(n4562), .O(n4563)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6765.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6766 (.I0(n3953), .I1(n3923), .I2(n4490), .I3(n4477), 
            .O(n4564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6766.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6767 (.I0(n4556), .I1(n4558), .I2(n4563), .I3(n4564), 
            .O(n3656)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6767.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6768 (.I0(n3933), .I1(n4221), .I2(n3920), .I3(n3921), 
            .O(n4565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6768.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6769 (.I0(n3945), .I1(n4412), .I2(n4450), .I3(n4565), 
            .O(n4566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__6769.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__6770 (.I0(n3943), .I1(n3945), .I2(n3917), .I3(n4428), 
            .O(n4567)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__6770.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__6771 (.I0(n4418), .I1(n4542), .I2(n4566), .I3(n4567), 
            .O(n3659)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6771.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6772 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[6] ), 
            .I2(\useone/round_flag[5] ), .O(n4568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6772.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6773 (.I0(n4568), .I1(n3901), .I2(\useone/round_flag[2] ), 
            .I3(\useone/round_flag[0] ), .O(n4569)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6773.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6774 (.I0(\useone/round_flag[3] ), .I1(n4298), .I2(n4228), 
            .I3(\useone/round_flag[2] ), .O(n4570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3dcf */ ;
    defparam LUT__6774.LUTMASK = 16'h3dcf;
    EFX_LUT4 LUT__6775 (.I0(n4459), .I1(n4570), .I2(n3926), .I3(n4539), 
            .O(n4571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6775.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6776 (.I0(\useone/round_flag[1] ), .I1(n4266), .I2(n3917), 
            .O(n4572)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6776.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6777 (.I0(n4440), .I1(n4572), .I2(n3953), .I3(n3903), 
            .O(n4573)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0ff1 */ ;
    defparam LUT__6777.LUTMASK = 16'h0ff1;
    EFX_LUT4 LUT__6778 (.I0(n3903), .I1(n3933), .I2(\useone/round_flag[0] ), 
            .I3(n3943), .O(n4574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6778.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6779 (.I0(n4574), .I1(n4532), .I2(n4533), .I3(n4438), 
            .O(n4575)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__6779.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__6780 (.I0(n4569), .I1(n4571), .I2(n4573), .I3(n4575), 
            .O(n3662)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6780.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6781 (.I0(n3917), .I1(\useone/round_flag[0] ), .I2(n3927), 
            .I3(\useone/round_flag[1] ), .O(n4576)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc83f */ ;
    defparam LUT__6781.LUTMASK = 16'hc83f;
    EFX_LUT4 LUT__6782 (.I0(n3918), .I1(\useone/round_flag[0] ), .O(n4577)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__6782.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__6783 (.I0(n4576), .I1(n4577), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[2] ), .O(n4578)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hadc0 */ ;
    defparam LUT__6783.LUTMASK = 16'hadc0;
    EFX_LUT4 LUT__6784 (.I0(\useone/round_flag[0] ), .I1(n3943), .I2(n3901), 
            .I3(n4508), .O(n4579)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__6784.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__6785 (.I0(n3918), .I1(n3924), .I2(\useone/round_flag[1] ), 
            .I3(n4510), .O(n4580)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hca00 */ ;
    defparam LUT__6785.LUTMASK = 16'hca00;
    EFX_LUT4 LUT__6786 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[1] ), 
            .I2(\useone/round_flag[4] ), .O(n4581)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6786.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6787 (.I0(\useone/round_flag[0] ), .I1(n3917), .I2(n4412), 
            .I3(n4581), .O(n4582)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6787.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6788 (.I0(n3913), .I1(n3933), .I2(n4582), .I3(n3938), 
            .O(n4583)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0700 */ ;
    defparam LUT__6788.LUTMASK = 16'h0700;
    EFX_LUT4 LUT__6789 (.I0(n4578), .I1(n4580), .I2(n4579), .I3(n4583), 
            .O(n3665)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefff */ ;
    defparam LUT__6789.LUTMASK = 16'hefff;
    EFX_LUT4 LUT__6790 (.I0(n3927), .I1(n4479), .I2(n3918), .I3(n3953), 
            .O(n4584)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6790.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6791 (.I0(n3903), .I1(n4479), .I2(n4440), .I3(n4584), 
            .O(n4585)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6791.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6792 (.I0(n4402), .I1(n3917), .I2(\useone/round_flag[0] ), 
            .I3(n3937), .O(n4586)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6792.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6793 (.I0(n4586), .I1(n3926), .I2(n4547), .O(n4587)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6793.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6794 (.I0(n3927), .I1(n3953), .I2(n3917), .I3(n3943), 
            .O(n4588)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6794.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6795 (.I0(n3903), .I1(n3914), .I2(n3918), .I3(n3913), 
            .O(n4589)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6795.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6796 (.I0(n4480), .I1(n4500), .I2(n4588), .I3(n4589), 
            .O(n4590)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__6796.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__6797 (.I0(n4585), .I1(n4587), .I2(n4590), .I3(n4417), 
            .O(n3668)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6797.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6798 (.I0(n3933), .I1(\useone/round_flag[1] ), .I2(n3918), 
            .I3(\useone/round_flag[2] ), .O(n4591)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__6798.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__6799 (.I0(n4591), .I1(\useone/round_flag[0] ), .O(n4592)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6799.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6800 (.I0(\useone/round_flag[2] ), .I1(n3923), .I2(n3909), 
            .O(n4593)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6800.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6801 (.I0(n3924), .I1(n3943), .I2(n4472), .I3(n4593), 
            .O(n4594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__6801.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__6802 (.I0(n3927), .I1(n3933), .I2(\useone/round_flag[1] ), 
            .O(n4595)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6802.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6803 (.I0(\useone/n46233 ), .I1(n3903), .I2(n4595), 
            .I3(\useone/round_flag[2] ), .O(n4596)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbf0 */ ;
    defparam LUT__6803.LUTMASK = 16'hbbf0;
    EFX_LUT4 LUT__6804 (.I0(\useone/round_flag[4] ), .I1(n4221), .I2(n3937), 
            .O(n4597)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6804.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6805 (.I0(n4402), .I1(n4597), .I2(n4462), .I3(n4588), 
            .O(n4598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d00 */ ;
    defparam LUT__6805.LUTMASK = 16'h0d00;
    EFX_LUT4 LUT__6806 (.I0(n4592), .I1(n4594), .I2(n4596), .I3(n4598), 
            .O(n3671)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6806.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6807 (.I0(n3901), .I1(\useone/round_flag[0] ), .I2(n3923), 
            .I3(\useone/round_flag[1] ), .O(n4599)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcf15 */ ;
    defparam LUT__6807.LUTMASK = 16'hcf15;
    EFX_LUT4 LUT__6808 (.I0(n3928), .I1(n3917), .I2(n4599), .I3(\useone/round_flag[2] ), 
            .O(n4600)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__6808.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__6809 (.I0(n3932), .I1(n3949), .I2(n3918), .O(n4601)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6809.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6810 (.I0(n3927), .I1(n3924), .I2(\useone/round_flag[2] ), 
            .I3(n3909), .O(n4602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0c0a */ ;
    defparam LUT__6810.LUTMASK = 16'h0c0a;
    EFX_LUT4 LUT__6811 (.I0(n3917), .I1(\useone/round_flag[2] ), .I2(n3927), 
            .I3(\useone/round_flag[0] ), .O(n4603)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__6811.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__6812 (.I0(n4413), .I1(n4601), .I2(n4602), .I3(n4603), 
            .O(n4604)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6812.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6813 (.I0(n4600), .I1(n4531), .I2(n4604), .I3(n3908), 
            .O(n3674)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6813.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6814 (.I0(n3933), .I1(n3918), .I2(\useone/round_flag[0] ), 
            .I3(n4254), .O(n4605)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6814.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6815 (.I0(\useone/round_flag[4] ), .I1(n3928), .I2(n4543), 
            .O(n4606)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__6815.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__6816 (.I0(n3933), .I1(n4221), .I2(n3937), .I3(n4402), 
            .O(n4607)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6816.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6817 (.I0(n3924), .I1(n3937), .I2(n4446), .I3(n4242), 
            .O(n4608)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6817.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6818 (.I0(n4605), .I1(n4606), .I2(n4607), .I3(n4608), 
            .O(n4609)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6818.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6819 (.I0(n4573), .I1(n4489), .I2(n4422), .I3(n4609), 
            .O(n3677)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6819.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6820 (.I0(\useone/round_flag[0] ), .I1(n3927), .I2(n3924), 
            .I3(\useone/round_flag[1] ), .O(n4610)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0f57 */ ;
    defparam LUT__6820.LUTMASK = 16'h0f57;
    EFX_LUT4 LUT__6821 (.I0(n3903), .I1(n3901), .I2(\useone/n46233 ), 
            .O(n4611)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6821.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6822 (.I0(n4611), .I1(n4610), .I2(\useone/round_flag[2] ), 
            .O(n4612)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__6822.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__6823 (.I0(n4511), .I1(n4549), .I2(n4589), .O(n4613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6823.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6824 (.I0(n4612), .I1(n4456), .I2(n4613), .I3(n4405), 
            .O(n3680)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6824.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6825 (.I0(n4574), .I1(n4438), .O(n4614)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6825.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6826 (.I0(n3943), .I1(n3932), .O(n4615)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__6826.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__6827 (.I0(n3953), .I1(n3945), .I2(n3923), .O(n4616)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6827.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6828 (.I0(n3912), .I1(n4615), .I2(n4616), .O(n4617)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__6828.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__6829 (.I0(\useone/round_flag[2] ), .I1(n3917), .I2(n3918), 
            .O(n4618)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6829.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6830 (.I0(\useone/round_flag[1] ), .I1(n3924), .I2(n4482), 
            .I3(n4618), .O(n4619)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7000 */ ;
    defparam LUT__6830.LUTMASK = 16'h7000;
    EFX_LUT4 LUT__6831 (.I0(n4242), .I1(n3905), .I2(\useone/round_flag[1] ), 
            .I3(n3917), .O(n4620)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7077 */ ;
    defparam LUT__6831.LUTMASK = 16'h7077;
    EFX_LUT4 LUT__6832 (.I0(n3902), .I1(n3903), .I2(n3925), .I3(n3924), 
            .O(n4621)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6832.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6833 (.I0(n4593), .I1(n4620), .I2(n4621), .O(n4622)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6833.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6834 (.I0(n4614), .I1(n4617), .I2(n4619), .I3(n4622), 
            .O(n3683)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6834.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6835 (.I0(n3933), .I1(n4266), .I2(\useone/round_flag[1] ), 
            .I3(n4221), .O(n4623)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'haf0c */ ;
    defparam LUT__6835.LUTMASK = 16'haf0c;
    EFX_LUT4 LUT__6836 (.I0(n3953), .I1(\useone/round_flag[1] ), .I2(n4623), 
            .I3(n3918), .O(n4624)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfac0 */ ;
    defparam LUT__6836.LUTMASK = 16'hfac0;
    EFX_LUT4 LUT__6837 (.I0(n3903), .I1(n3933), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[0] ), .O(n4625)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6837.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6838 (.I0(n4266), .I1(n4254), .I2(n3901), .O(n4626)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6838.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6839 (.I0(n3923), .I1(n3917), .I2(n3937), .O(n4627)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__6839.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__6840 (.I0(n4625), .I1(n4626), .I2(n4453), .I3(n4627), 
            .O(n4628)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6840.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6841 (.I0(\useone/n46233 ), .I1(n3903), .I2(\useone/round_flag[2] ), 
            .I3(n4499), .O(n4629)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__6841.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__6842 (.I0(n4624), .I1(n4628), .I2(n4552), .I3(n4629), 
            .O(n3686)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6842.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6843 (.I0(\useone/round_flag[1] ), .I1(\useone/round_flag[2] ), 
            .I2(\useone/round_flag[4] ), .I3(\useone/round_flag[5] ), .O(n4630)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5b3c */ ;
    defparam LUT__6843.LUTMASK = 16'h5b3c;
    EFX_LUT4 LUT__6844 (.I0(n4630), .I1(\useone/round_flag[0] ), .I2(n4559), 
            .O(n4631)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6844.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6845 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[2] ), .I3(\useone/round_flag[4] ), .O(n4632)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbecf */ ;
    defparam LUT__6845.LUTMASK = 16'hbecf;
    EFX_LUT4 LUT__6846 (.I0(n4632), .I1(\useone/round_flag[1] ), .I2(n4459), 
            .O(n4633)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__6846.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__6847 (.I0(n4494), .I1(n4515), .I2(n4605), .I3(n4633), 
            .O(n4634)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__6847.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__6848 (.I0(n4631), .I1(n4617), .I2(n4634), .I3(n4596), 
            .O(n3689)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbfff */ ;
    defparam LUT__6848.LUTMASK = 16'hbfff;
    EFX_LUT4 LUT__6849 (.I0(n3901), .I1(n3923), .I2(n3927), .I3(\useone/round_flag[2] ), 
            .O(n4635)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0305 */ ;
    defparam LUT__6849.LUTMASK = 16'h0305;
    EFX_LUT4 LUT__6850 (.I0(n3905), .I1(n4254), .I2(n3925), .O(n4636)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0707 */ ;
    defparam LUT__6850.LUTMASK = 16'h0707;
    EFX_LUT4 LUT__6851 (.I0(\useone/round_flag[0] ), .I1(n4635), .I2(n4636), 
            .O(n4637)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__6851.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__6852 (.I0(\useone/round_flag[2] ), .I1(\useone/round_flag[4] ), 
            .I2(n3909), .I3(n4402), .O(n4638)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6000 */ ;
    defparam LUT__6852.LUTMASK = 16'h6000;
    EFX_LUT4 LUT__6853 (.I0(n4526), .I1(n3924), .O(n4639)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6853.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6854 (.I0(\useone/round_flag[2] ), .I1(n4402), .I2(n3903), 
            .I3(n3928), .O(n4640)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__6854.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__6855 (.I0(n3909), .I1(n3903), .I2(n3917), .I3(n4266), 
            .O(n4641)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6855.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6856 (.I0(n4639), .I1(n4640), .I2(n4641), .I3(n4620), 
            .O(n4642)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__6856.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__6857 (.I0(\useone/round_flag[0] ), .I1(\useone/round_flag[3] ), 
            .I2(\useone/round_flag[1] ), .I3(\useone/round_flag[2] ), .O(n4643)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0110 */ ;
    defparam LUT__6857.LUTMASK = 16'h0110;
    EFX_LUT4 LUT__6858 (.I0(n3912), .I1(n4643), .I2(n3933), .I3(n4503), 
            .O(n4644)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0777 */ ;
    defparam LUT__6858.LUTMASK = 16'h0777;
    EFX_LUT4 LUT__6859 (.I0(n4637), .I1(n4638), .I2(n4642), .I3(n4644), 
            .O(n3692)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefff */ ;
    defparam LUT__6859.LUTMASK = 16'hefff;
    EFX_LUT4 LUT__6860 (.I0(n3917), .I1(n3902), .I2(n3933), .I3(\useone/round_flag[0] ), 
            .O(n4645)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00f8 */ ;
    defparam LUT__6860.LUTMASK = 16'h00f8;
    EFX_LUT4 LUT__6861 (.I0(n4645), .I1(n4467), .I2(n4441), .O(n4646)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__6861.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__6862 (.I0(n4527), .I1(n3900), .I2(n3924), .O(n4647)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__6862.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__6863 (.I0(n3933), .I1(n3917), .I2(\useone/round_flag[1] ), 
            .I3(\useone/round_flag[2] ), .O(n4648)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ff3 */ ;
    defparam LUT__6863.LUTMASK = 16'h5ff3;
    EFX_LUT4 LUT__6864 (.I0(n4577), .I1(n4626), .I2(n4647), .I3(n4648), 
            .O(n4649)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6864.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6865 (.I0(n4487), .I1(n4583), .I2(n4646), .I3(n4649), 
            .O(n3695)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6865.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6866 (.I0(n3937), .I1(n3917), .O(n4650)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__6866.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__6867 (.I0(n3924), .I1(n3933), .I2(\useone/round_flag[2] ), 
            .I3(n3931), .O(n4651)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac00 */ ;
    defparam LUT__6867.LUTMASK = 16'hac00;
    EFX_LUT4 LUT__6868 (.I0(n4455), .I1(n4650), .I2(n4651), .I3(n4644), 
            .O(n4652)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__6868.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__6869 (.I0(n3918), .I1(n4615), .I2(n4504), .I3(n4486), 
            .O(n4653)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h000d */ ;
    defparam LUT__6869.LUTMASK = 16'h000d;
    EFX_LUT4 LUT__6870 (.I0(n4594), .I1(n4652), .I2(n4653), .I3(n4529), 
            .O(n3698)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__6870.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__6871 (.I0(\useone/g[31] ), .I1(\useone/f[31] ), .I2(\useone/e[31] ), 
            .O(n3701)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6871.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6872 (.I0(\useone/f[30] ), .I1(\useone/g[30] ), .I2(\useone/e[30] ), 
            .O(n3704)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6872.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6873 (.I0(\useone/g[29] ), .I1(\useone/f[29] ), .I2(\useone/e[29] ), 
            .O(n3707)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6873.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6874 (.I0(\useone/f[28] ), .I1(\useone/g[28] ), .I2(\useone/e[28] ), 
            .O(n3710)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6874.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6875 (.I0(\useone/g[27] ), .I1(\useone/f[27] ), .I2(\useone/e[27] ), 
            .O(n3713)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6875.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6876 (.I0(\useone/g[26] ), .I1(\useone/f[26] ), .I2(\useone/e[26] ), 
            .O(n3716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6876.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6877 (.I0(\useone/g[25] ), .I1(\useone/f[25] ), .I2(\useone/e[25] ), 
            .O(n3719)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6877.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6878 (.I0(\useone/f[24] ), .I1(\useone/g[24] ), .I2(\useone/e[24] ), 
            .O(n3722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6878.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6879 (.I0(\useone/g[23] ), .I1(\useone/f[23] ), .I2(\useone/e[23] ), 
            .O(n3725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6879.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6880 (.I0(\useone/g[22] ), .I1(\useone/f[22] ), .I2(\useone/e[22] ), 
            .O(n3728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6880.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6881 (.I0(\useone/g[21] ), .I1(\useone/f[21] ), .I2(\useone/e[21] ), 
            .O(n3731)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6881.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6882 (.I0(\useone/g[20] ), .I1(\useone/f[20] ), .I2(\useone/e[20] ), 
            .O(n3734)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6882.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6883 (.I0(\useone/f[19] ), .I1(\useone/g[19] ), .I2(\useone/e[19] ), 
            .O(n3737)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6883.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6884 (.I0(\useone/f[18] ), .I1(\useone/g[18] ), .I2(\useone/e[18] ), 
            .O(n3740)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6884.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6885 (.I0(\useone/f[17] ), .I1(\useone/g[17] ), .I2(\useone/e[17] ), 
            .O(n3743)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6885.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6886 (.I0(\useone/g[16] ), .I1(\useone/f[16] ), .I2(\useone/e[16] ), 
            .O(n3746)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6886.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6887 (.I0(\useone/g[15] ), .I1(\useone/f[15] ), .I2(\useone/e[15] ), 
            .O(n3749)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6887.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6888 (.I0(\useone/f[14] ), .I1(\useone/g[14] ), .I2(\useone/e[14] ), 
            .O(n3752)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6888.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6889 (.I0(\useone/g[13] ), .I1(\useone/f[13] ), .I2(\useone/e[13] ), 
            .O(n3755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6889.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6890 (.I0(\useone/f[12] ), .I1(\useone/g[12] ), .I2(\useone/e[12] ), 
            .O(n3758)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6890.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6891 (.I0(\useone/g[11] ), .I1(\useone/f[11] ), .I2(\useone/e[11] ), 
            .O(n3761)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6891.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6892 (.I0(\useone/g[10] ), .I1(\useone/f[10] ), .I2(\useone/e[10] ), 
            .O(n3764)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6892.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6893 (.I0(\useone/f[9] ), .I1(\useone/g[9] ), .I2(\useone/e[9] ), 
            .O(n3767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6893.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6894 (.I0(\useone/g[8] ), .I1(\useone/f[8] ), .I2(\useone/e[8] ), 
            .O(n3770)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6894.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6895 (.I0(\useone/g[7] ), .I1(\useone/f[7] ), .I2(\useone/e[7] ), 
            .O(n3773)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6895.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6896 (.I0(\useone/f[6] ), .I1(\useone/g[6] ), .I2(\useone/e[6] ), 
            .O(n3776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6896.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6897 (.I0(\useone/f[5] ), .I1(\useone/g[5] ), .I2(\useone/e[5] ), 
            .O(n3779)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6897.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6898 (.I0(\useone/f[4] ), .I1(\useone/g[4] ), .I2(\useone/e[4] ), 
            .O(n3782)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__6898.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__6899 (.I0(\useone/f[3] ), .I1(\useone/g[3] ), .I2(\useone/e[3] ), 
            .O(n3785)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__6899.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__6900 (.I0(\useone/f[2] ), .I1(\useone/g[2] ), .I2(\useone/e[2] ), 
            .O(n3788)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hc5c5 */ ;
    defparam LUT__6900.LUTMASK = 16'hc5c5;
    EFX_LUT4 LUT__6901 (.I0(\useone/f[1] ), .I1(\useone/g[1] ), .I2(\useone/e[1] ), 
            .O(n3791)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3a3a */ ;
    defparam LUT__6901.LUTMASK = 16'h3a3a;
    EFX_LUT4 LUT__6902 (.I0(\useone/e[5] ), .I1(\useone/e[10] ), .I2(\useone/e[24] ), 
            .O(n3793)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6902.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6903 (.I0(\useone/e[4] ), .I1(\useone/e[9] ), .I2(\useone/e[23] ), 
            .O(n3795)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6903.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6904 (.I0(\useone/e[3] ), .I1(\useone/e[8] ), .I2(\useone/e[22] ), 
            .O(n3797)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6904.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6905 (.I0(\useone/e[2] ), .I1(\useone/e[7] ), .I2(\useone/e[21] ), 
            .O(n3799)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6905.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6906 (.I0(\useone/e[1] ), .I1(\useone/e[6] ), .I2(\useone/e[20] ), 
            .O(n3801)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6906.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6907 (.I0(\useone/e[0] ), .I1(\useone/e[5] ), .I2(\useone/e[19] ), 
            .O(n3803)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6907.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6908 (.I0(\useone/e[4] ), .I1(\useone/e[18] ), .I2(\useone/e[31] ), 
            .O(n3805)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6908.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6909 (.I0(\useone/e[3] ), .I1(\useone/e[17] ), .I2(\useone/e[30] ), 
            .O(n3807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6909.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6910 (.I0(\useone/e[2] ), .I1(\useone/e[16] ), .I2(\useone/e[29] ), 
            .O(n3809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6910.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6911 (.I0(\useone/e[1] ), .I1(\useone/e[15] ), .I2(\useone/e[28] ), 
            .O(n3811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6911.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6912 (.I0(\useone/e[0] ), .I1(\useone/e[14] ), .I2(\useone/e[27] ), 
            .O(n3813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6912.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6913 (.I0(\useone/e[13] ), .I1(\useone/e[26] ), .I2(\useone/e[31] ), 
            .O(n3815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6913.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6914 (.I0(\useone/e[12] ), .I1(\useone/e[25] ), .I2(\useone/e[30] ), 
            .O(n3817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6914.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6915 (.I0(\useone/e[11] ), .I1(\useone/e[24] ), .I2(\useone/e[29] ), 
            .O(n3819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6915.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6916 (.I0(\useone/e[10] ), .I1(\useone/e[23] ), .I2(\useone/e[28] ), 
            .O(n3821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6916.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6917 (.I0(\useone/e[9] ), .I1(\useone/e[22] ), .I2(\useone/e[27] ), 
            .O(n3823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6917.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6918 (.I0(\useone/e[8] ), .I1(\useone/e[21] ), .I2(\useone/e[26] ), 
            .O(n3825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6918.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6919 (.I0(\useone/e[7] ), .I1(\useone/e[20] ), .I2(\useone/e[25] ), 
            .O(n3827)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6919.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6920 (.I0(\useone/e[6] ), .I1(\useone/e[19] ), .I2(\useone/e[24] ), 
            .O(n3829)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6920.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6921 (.I0(\useone/e[5] ), .I1(\useone/e[18] ), .I2(\useone/e[23] ), 
            .O(n3831)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6921.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6922 (.I0(\useone/e[4] ), .I1(\useone/e[17] ), .I2(\useone/e[22] ), 
            .O(n3833)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6922.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6923 (.I0(\useone/e[3] ), .I1(\useone/e[16] ), .I2(\useone/e[21] ), 
            .O(n3835)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6923.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6924 (.I0(\useone/e[2] ), .I1(\useone/e[15] ), .I2(\useone/e[20] ), 
            .O(n3837)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6924.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6925 (.I0(\useone/e[1] ), .I1(\useone/e[14] ), .I2(\useone/e[19] ), 
            .O(n3839)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6925.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6926 (.I0(\useone/e[0] ), .I1(\useone/e[13] ), .I2(\useone/e[18] ), 
            .O(n3841)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6926.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6927 (.I0(\useone/e[12] ), .I1(\useone/e[17] ), .I2(\useone/e[31] ), 
            .O(n3843)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6927.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6928 (.I0(\useone/e[11] ), .I1(\useone/e[16] ), .I2(\useone/e[30] ), 
            .O(n3845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6928.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6929 (.I0(\useone/e[10] ), .I1(\useone/e[15] ), .I2(\useone/e[29] ), 
            .O(n3847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6929.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6930 (.I0(\useone/e[9] ), .I1(\useone/e[14] ), .I2(\useone/e[28] ), 
            .O(n3849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6930.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6931 (.I0(\useone/e[8] ), .I1(\useone/e[13] ), .I2(\useone/e[27] ), 
            .O(n3851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__6931.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__6932 (.I0(\useone/e[7] ), .I1(\useone/e[12] ), .I2(\useone/e[26] ), 
            .O(n3853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6969 */ ;
    defparam LUT__6932.LUTMASK = 16'h6969;
    EFX_LUT4 LUT__6935 (.I0(o_uart_tx_2), .O(o_uart_tx)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__6935.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__5631 (.I0(o_Tx_active), .I1(\state[1] ), .I2(\state[0] ), 
            .O(ceg_net40)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__5631.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__5632 (.I0(\state[0] ), .I1(\state[1] ), .O(ceg_net85)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__5632.LUTMASK = 16'h8888;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(clk), .O(\clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_FF_d7ffea96_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_d7ffea96_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_d7ffea96_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_d7ffea96_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_d7ffea96_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_d7ffea96_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_d7ffea96_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_d7ffea96_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_d7ffea96_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_d7ffea96_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_d7ffea96_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_221
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_222
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_223
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_224
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_225
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_226
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_227
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_228
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_229
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_230
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_231
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_232
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_233
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_234
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_235
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_d7ffea96_236
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_d7ffea96_0
// module not written out since it is a black box. 
//

